module VCR( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output        io_host_aw_ready, // @[:@6.4]
  input         io_host_aw_valid, // @[:@6.4]
  input  [15:0] io_host_aw_bits_addr, // @[:@6.4]
  output        io_host_w_ready, // @[:@6.4]
  input         io_host_w_valid, // @[:@6.4]
  input  [31:0] io_host_w_bits_data, // @[:@6.4]
  input         io_host_b_ready, // @[:@6.4]
  output        io_host_b_valid, // @[:@6.4]
  output        io_host_ar_ready, // @[:@6.4]
  input         io_host_ar_valid, // @[:@6.4]
  input  [15:0] io_host_ar_bits_addr, // @[:@6.4]
  input         io_host_r_ready, // @[:@6.4]
  output        io_host_r_valid, // @[:@6.4]
  output [31:0] io_host_r_bits_data, // @[:@6.4]
  output        io_vcr_launch, // @[:@6.4]
  input         io_vcr_finish, // @[:@6.4]
  input         io_vcr_ecnt_0_valid, // @[:@6.4]
  input  [31:0] io_vcr_ecnt_0_bits, // @[:@6.4]
  output [31:0] io_vcr_vals_0, // @[:@6.4]
  output [31:0] io_vcr_ptrs_0, // @[:@6.4]
  output [31:0] io_vcr_ptrs_1, // @[:@6.4]
  output [31:0] io_vcr_ptrs_2, // @[:@6.4]
  output [31:0] io_vcr_ptrs_3, // @[:@6.4]
  output [31:0] io_vcr_ptrs_4, // @[:@6.4]
  output [31:0] io_vcr_ptrs_5, // @[:@6.4]
  input         io_vcr_ucnt_0_valid, // @[:@6.4]
  input  [31:0] io_vcr_ucnt_0_bits // @[:@6.4]
);
  reg [15:0] waddr; // @[VCR.scala 94:22:@8.4]
  reg [31:0] _RAND_0;
  reg [1:0] wstate; // @[VCR.scala 97:23:@9.4]
  reg [31:0] _RAND_1;
  reg  rstate; // @[VCR.scala 101:23:@10.4]
  reg [31:0] _RAND_2;
  reg [31:0] rdata; // @[VCR.scala 102:22:@11.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_0; // @[VCR.scala 108:37:@12.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_1; // @[VCR.scala 108:37:@13.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_2; // @[VCR.scala 108:37:@14.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_3; // @[VCR.scala 108:37:@15.4]
  reg [31:0] _RAND_7;
  reg [31:0] reg_4; // @[VCR.scala 108:37:@16.4]
  reg [31:0] _RAND_8;
  reg [31:0] reg_5; // @[VCR.scala 108:37:@17.4]
  reg [31:0] _RAND_9;
  reg [31:0] reg_6; // @[VCR.scala 108:37:@18.4]
  reg [31:0] _RAND_10;
  reg [31:0] reg_7; // @[VCR.scala 108:37:@19.4]
  reg [31:0] _RAND_11;
  reg [31:0] reg_8; // @[VCR.scala 108:37:@20.4]
  reg [31:0] _RAND_12;
  reg [31:0] reg_9; // @[VCR.scala 108:37:@21.4]
  reg [31:0] _RAND_13;
  wire  _T_159; // @[Conditional.scala 37:30:@22.4]
  wire [1:0] _GEN_0; // @[VCR.scala 118:30:@24.6]
  wire  _T_160; // @[Conditional.scala 37:30:@29.6]
  wire [1:0] _GEN_1; // @[VCR.scala 123:29:@31.8]
  wire  _T_161; // @[Conditional.scala 37:30:@36.8]
  wire [1:0] _GEN_2; // @[VCR.scala 128:29:@38.10]
  wire [1:0] _GEN_3; // @[Conditional.scala 39:67:@37.8]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@30.6]
  wire [1:0] _GEN_5; // @[Conditional.scala 40:58:@23.4]
  wire  _T_162; // @[Decoupled.scala 37:37:@42.4]
  wire [15:0] _GEN_6; // @[VCR.scala 134:27:@43.4]
  wire  _T_167; // @[Conditional.scala 37:30:@53.4]
  wire  _GEN_7; // @[VCR.scala 143:30:@55.6]
  wire  _GEN_8; // @[VCR.scala 148:29:@62.8]
  wire  _GEN_9; // @[Conditional.scala 39:67:@61.6]
  wire  _GEN_10; // @[Conditional.scala 40:58:@54.4]
  wire  _T_173; // @[Decoupled.scala 37:37:@76.6]
  wire  _T_175; // @[VCR.scala 161:44:@77.6]
  wire  _T_176; // @[VCR.scala 161:31:@78.6]
  wire [31:0] _GEN_11; // @[VCR.scala 161:55:@79.6]
  wire [31:0] _GEN_12; // @[VCR.scala 159:23:@72.4]
  wire  _T_179; // @[VCR.scala 168:51:@87.6]
  wire  _T_180; // @[VCR.scala 168:33:@88.6]
  wire [31:0] _GEN_13; // @[VCR.scala 168:62:@89.6]
  wire [31:0] _GEN_14; // @[VCR.scala 166:32:@82.4]
  wire  _T_183; // @[VCR.scala 174:45:@93.4]
  wire  _T_184; // @[VCR.scala 174:27:@94.4]
  wire [31:0] _GEN_15; // @[VCR.scala 174:56:@95.4]
  wire  _T_187; // @[VCR.scala 174:45:@99.4]
  wire  _T_188; // @[VCR.scala 174:27:@100.4]
  wire [31:0] _GEN_16; // @[VCR.scala 174:56:@101.4]
  wire  _T_191; // @[VCR.scala 174:45:@105.4]
  wire  _T_192; // @[VCR.scala 174:27:@106.4]
  wire [31:0] _GEN_17; // @[VCR.scala 174:56:@107.4]
  wire  _T_195; // @[VCR.scala 174:45:@111.4]
  wire  _T_196; // @[VCR.scala 174:27:@112.4]
  wire [31:0] _GEN_18; // @[VCR.scala 174:56:@113.4]
  wire  _T_199; // @[VCR.scala 174:45:@117.4]
  wire  _T_200; // @[VCR.scala 174:27:@118.4]
  wire [31:0] _GEN_19; // @[VCR.scala 174:56:@119.4]
  wire  _T_203; // @[VCR.scala 174:45:@123.4]
  wire  _T_204; // @[VCR.scala 174:27:@124.4]
  wire [31:0] _GEN_20; // @[VCR.scala 174:56:@125.4]
  wire  _T_207; // @[VCR.scala 174:45:@129.4]
  wire  _T_208; // @[VCR.scala 174:27:@130.4]
  wire [31:0] _GEN_21; // @[VCR.scala 174:56:@131.4]
  wire  _T_209; // @[Decoupled.scala 37:37:@134.4]
  wire  _T_211; // @[Mux.scala 46:19:@136.6]
  wire [31:0] _T_212; // @[Mux.scala 46:16:@137.6]
  wire  _T_213; // @[Mux.scala 46:19:@138.6]
  wire [31:0] _T_214; // @[Mux.scala 46:16:@139.6]
  wire  _T_215; // @[Mux.scala 46:19:@140.6]
  wire [31:0] _T_216; // @[Mux.scala 46:16:@141.6]
  wire  _T_217; // @[Mux.scala 46:19:@142.6]
  wire [31:0] _T_218; // @[Mux.scala 46:16:@143.6]
  wire  _T_219; // @[Mux.scala 46:19:@144.6]
  wire [31:0] _T_220; // @[Mux.scala 46:16:@145.6]
  wire  _T_221; // @[Mux.scala 46:19:@146.6]
  wire [31:0] _T_222; // @[Mux.scala 46:16:@147.6]
  wire  _T_223; // @[Mux.scala 46:19:@148.6]
  wire [31:0] _T_224; // @[Mux.scala 46:16:@149.6]
  wire  _T_225; // @[Mux.scala 46:19:@150.6]
  wire [31:0] _T_226; // @[Mux.scala 46:16:@151.6]
  wire  _T_227; // @[Mux.scala 46:19:@152.6]
  wire [31:0] _T_228; // @[Mux.scala 46:16:@153.6]
  wire  _T_229; // @[Mux.scala 46:19:@154.6]
  wire [31:0] _T_230; // @[Mux.scala 46:16:@155.6]
  wire [31:0] _GEN_22; // @[VCR.scala 179:27:@135.4]
  wire  _T_234; // @[VCR.scala 202:51:@172.6]
  wire  _T_235; // @[VCR.scala 202:33:@173.6]
  wire [31:0] _GEN_23; // @[VCR.scala 202:62:@174.6]
  wire [31:0] _GEN_24; // @[VCR.scala 200:32:@167.4]
  assign _T_159 = 2'h0 == wstate; // @[Conditional.scala 37:30:@22.4]
  assign _GEN_0 = io_host_aw_valid ? 2'h1 : wstate; // @[VCR.scala 118:30:@24.6]
  assign _T_160 = 2'h1 == wstate; // @[Conditional.scala 37:30:@29.6]
  assign _GEN_1 = io_host_w_valid ? 2'h2 : wstate; // @[VCR.scala 123:29:@31.8]
  assign _T_161 = 2'h2 == wstate; // @[Conditional.scala 37:30:@36.8]
  assign _GEN_2 = io_host_b_ready ? 2'h0 : wstate; // @[VCR.scala 128:29:@38.10]
  assign _GEN_3 = _T_161 ? _GEN_2 : wstate; // @[Conditional.scala 39:67:@37.8]
  assign _GEN_4 = _T_160 ? _GEN_1 : _GEN_3; // @[Conditional.scala 39:67:@30.6]
  assign _GEN_5 = _T_159 ? _GEN_0 : _GEN_4; // @[Conditional.scala 40:58:@23.4]
  assign _T_162 = io_host_aw_ready & io_host_aw_valid; // @[Decoupled.scala 37:37:@42.4]
  assign _GEN_6 = _T_162 ? io_host_aw_bits_addr : waddr; // @[VCR.scala 134:27:@43.4]
  assign _T_167 = 1'h0 == rstate; // @[Conditional.scala 37:30:@53.4]
  assign _GEN_7 = io_host_ar_valid ? 1'h1 : rstate; // @[VCR.scala 143:30:@55.6]
  assign _GEN_8 = io_host_r_ready ? 1'h0 : rstate; // @[VCR.scala 148:29:@62.8]
  assign _GEN_9 = rstate ? _GEN_8 : rstate; // @[Conditional.scala 39:67:@61.6]
  assign _GEN_10 = _T_167 ? _GEN_7 : _GEN_9; // @[Conditional.scala 40:58:@54.4]
  assign _T_173 = io_host_w_ready & io_host_w_valid; // @[Decoupled.scala 37:37:@76.6]
  assign _T_175 = 16'h0 == waddr; // @[VCR.scala 161:44:@77.6]
  assign _T_176 = _T_173 & _T_175; // @[VCR.scala 161:31:@78.6]
  assign _GEN_11 = _T_176 ? io_host_w_bits_data : reg_0; // @[VCR.scala 161:55:@79.6]
  assign _GEN_12 = io_vcr_finish ? 32'h2 : _GEN_11; // @[VCR.scala 159:23:@72.4]
  assign _T_179 = 16'h4 == waddr; // @[VCR.scala 168:51:@87.6]
  assign _T_180 = _T_173 & _T_179; // @[VCR.scala 168:33:@88.6]
  assign _GEN_13 = _T_180 ? io_host_w_bits_data : reg_1; // @[VCR.scala 168:62:@89.6]
  assign _GEN_14 = io_vcr_ecnt_0_valid ? io_vcr_ecnt_0_bits : _GEN_13; // @[VCR.scala 166:32:@82.4]
  assign _T_183 = 16'h8 == waddr; // @[VCR.scala 174:45:@93.4]
  assign _T_184 = _T_173 & _T_183; // @[VCR.scala 174:27:@94.4]
  assign _GEN_15 = _T_184 ? io_host_w_bits_data : reg_2; // @[VCR.scala 174:56:@95.4]
  assign _T_187 = 16'hc == waddr; // @[VCR.scala 174:45:@99.4]
  assign _T_188 = _T_173 & _T_187; // @[VCR.scala 174:27:@100.4]
  assign _GEN_16 = _T_188 ? io_host_w_bits_data : reg_3; // @[VCR.scala 174:56:@101.4]
  assign _T_191 = 16'h10 == waddr; // @[VCR.scala 174:45:@105.4]
  assign _T_192 = _T_173 & _T_191; // @[VCR.scala 174:27:@106.4]
  assign _GEN_17 = _T_192 ? io_host_w_bits_data : reg_4; // @[VCR.scala 174:56:@107.4]
  assign _T_195 = 16'h14 == waddr; // @[VCR.scala 174:45:@111.4]
  assign _T_196 = _T_173 & _T_195; // @[VCR.scala 174:27:@112.4]
  assign _GEN_18 = _T_196 ? io_host_w_bits_data : reg_5; // @[VCR.scala 174:56:@113.4]
  assign _T_199 = 16'h18 == waddr; // @[VCR.scala 174:45:@117.4]
  assign _T_200 = _T_173 & _T_199; // @[VCR.scala 174:27:@118.4]
  assign _GEN_19 = _T_200 ? io_host_w_bits_data : reg_6; // @[VCR.scala 174:56:@119.4]
  assign _T_203 = 16'h1c == waddr; // @[VCR.scala 174:45:@123.4]
  assign _T_204 = _T_173 & _T_203; // @[VCR.scala 174:27:@124.4]
  assign _GEN_20 = _T_204 ? io_host_w_bits_data : reg_7; // @[VCR.scala 174:56:@125.4]
  assign _T_207 = 16'h20 == waddr; // @[VCR.scala 174:45:@129.4]
  assign _T_208 = _T_173 & _T_207; // @[VCR.scala 174:27:@130.4]
  assign _GEN_21 = _T_208 ? io_host_w_bits_data : reg_8; // @[VCR.scala 174:56:@131.4]
  assign _T_209 = io_host_ar_ready & io_host_ar_valid; // @[Decoupled.scala 37:37:@134.4]
  assign _T_211 = 16'h24 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@136.6]
  assign _T_212 = _T_211 ? reg_9 : 32'h0; // @[Mux.scala 46:16:@137.6]
  assign _T_213 = 16'h20 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@138.6]
  assign _T_214 = _T_213 ? reg_8 : _T_212; // @[Mux.scala 46:16:@139.6]
  assign _T_215 = 16'h1c == io_host_ar_bits_addr; // @[Mux.scala 46:19:@140.6]
  assign _T_216 = _T_215 ? reg_7 : _T_214; // @[Mux.scala 46:16:@141.6]
  assign _T_217 = 16'h18 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@142.6]
  assign _T_218 = _T_217 ? reg_6 : _T_216; // @[Mux.scala 46:16:@143.6]
  assign _T_219 = 16'h14 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@144.6]
  assign _T_220 = _T_219 ? reg_5 : _T_218; // @[Mux.scala 46:16:@145.6]
  assign _T_221 = 16'h10 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@146.6]
  assign _T_222 = _T_221 ? reg_4 : _T_220; // @[Mux.scala 46:16:@147.6]
  assign _T_223 = 16'hc == io_host_ar_bits_addr; // @[Mux.scala 46:19:@148.6]
  assign _T_224 = _T_223 ? reg_3 : _T_222; // @[Mux.scala 46:16:@149.6]
  assign _T_225 = 16'h8 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@150.6]
  assign _T_226 = _T_225 ? reg_2 : _T_224; // @[Mux.scala 46:16:@151.6]
  assign _T_227 = 16'h4 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@152.6]
  assign _T_228 = _T_227 ? reg_1 : _T_226; // @[Mux.scala 46:16:@153.6]
  assign _T_229 = 16'h0 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@154.6]
  assign _T_230 = _T_229 ? reg_0 : _T_228; // @[Mux.scala 46:16:@155.6]
  assign _GEN_22 = _T_209 ? _T_230 : rdata; // @[VCR.scala 179:27:@135.4]
  assign _T_234 = 16'h24 == waddr; // @[VCR.scala 202:51:@172.6]
  assign _T_235 = _T_173 & _T_234; // @[VCR.scala 202:33:@173.6]
  assign _GEN_23 = _T_235 ? io_host_w_bits_data : reg_9; // @[VCR.scala 202:62:@174.6]
  assign _GEN_24 = io_vcr_ucnt_0_valid ? io_vcr_ucnt_0_bits : _GEN_23; // @[VCR.scala 200:32:@167.4]
  assign io_host_aw_ready = wstate == 2'h0; // @[VCR.scala 136:20:@47.4]
  assign io_host_w_ready = wstate == 2'h1; // @[VCR.scala 137:19:@49.4]
  assign io_host_b_valid = wstate == 2'h2; // @[VCR.scala 138:19:@51.4]
  assign io_host_ar_ready = rstate == 1'h0; // @[VCR.scala 154:20:@67.4]
  assign io_host_r_valid = rstate; // @[VCR.scala 155:19:@69.4]
  assign io_host_r_bits_data = rdata; // @[VCR.scala 156:23:@70.4]
  assign io_vcr_launch = reg_0[0]; // @[VCR.scala 183:17:@159.4]
  assign io_vcr_vals_0 = reg_2; // @[VCR.scala 186:20:@160.4]
  assign io_vcr_ptrs_0 = reg_3; // @[VCR.scala 191:22:@161.4]
  assign io_vcr_ptrs_1 = reg_4; // @[VCR.scala 191:22:@162.4]
  assign io_vcr_ptrs_2 = reg_5; // @[VCR.scala 191:22:@163.4]
  assign io_vcr_ptrs_3 = reg_6; // @[VCR.scala 191:22:@164.4]
  assign io_vcr_ptrs_4 = reg_7; // @[VCR.scala 191:22:@165.4]
  assign io_vcr_ptrs_5 = reg_8; // @[VCR.scala 191:22:@166.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waddr = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  wstate = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rstate = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  rdata = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_0 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_1 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_2 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_3 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_4 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_5 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_6 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_7 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  reg_8 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  reg_9 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      waddr <= 16'hffff;
    end else begin
      if (_T_162) begin
        waddr <= io_host_aw_bits_addr;
      end
    end
    if (reset) begin
      wstate <= 2'h0;
    end else begin
      if (_T_159) begin
        if (io_host_aw_valid) begin
          wstate <= 2'h1;
        end
      end else begin
        if (_T_160) begin
          if (io_host_w_valid) begin
            wstate <= 2'h2;
          end
        end else begin
          if (_T_161) begin
            if (io_host_b_ready) begin
              wstate <= 2'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      rstate <= 1'h0;
    end else begin
      if (_T_167) begin
        if (io_host_ar_valid) begin
          rstate <= 1'h1;
        end
      end else begin
        if (rstate) begin
          if (io_host_r_ready) begin
            rstate <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      rdata <= 32'h0;
    end else begin
      if (_T_209) begin
        if (_T_229) begin
          rdata <= reg_0;
        end else begin
          if (_T_227) begin
            rdata <= reg_1;
          end else begin
            if (_T_225) begin
              rdata <= reg_2;
            end else begin
              if (_T_223) begin
                rdata <= reg_3;
              end else begin
                if (_T_221) begin
                  rdata <= reg_4;
                end else begin
                  if (_T_219) begin
                    rdata <= reg_5;
                  end else begin
                    if (_T_217) begin
                      rdata <= reg_6;
                    end else begin
                      if (_T_215) begin
                        rdata <= reg_7;
                      end else begin
                        if (_T_213) begin
                          rdata <= reg_8;
                        end else begin
                          if (_T_211) begin
                            rdata <= reg_9;
                          end else begin
                            rdata <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_0 <= 32'h0;
    end else begin
      if (io_vcr_finish) begin
        reg_0 <= 32'h2;
      end else begin
        if (_T_176) begin
          reg_0 <= io_host_w_bits_data;
        end
      end
    end
    if (reset) begin
      reg_1 <= 32'h0;
    end else begin
      if (io_vcr_ecnt_0_valid) begin
        reg_1 <= io_vcr_ecnt_0_bits;
      end else begin
        if (_T_180) begin
          reg_1 <= io_host_w_bits_data;
        end
      end
    end
    if (reset) begin
      reg_2 <= 32'h0;
    end else begin
      if (_T_184) begin
        reg_2 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_3 <= 32'h0;
    end else begin
      if (_T_188) begin
        reg_3 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_4 <= 32'h0;
    end else begin
      if (_T_192) begin
        reg_4 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_5 <= 32'h0;
    end else begin
      if (_T_196) begin
        reg_5 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_6 <= 32'h0;
    end else begin
      if (_T_200) begin
        reg_6 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_7 <= 32'h0;
    end else begin
      if (_T_204) begin
        reg_7 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_8 <= 32'h0;
    end else begin
      if (_T_208) begin
        reg_8 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_9 <= 32'h0;
    end else begin
      if (io_vcr_ucnt_0_valid) begin
        reg_9 <= io_vcr_ucnt_0_bits;
      end else begin
        if (_T_235) begin
          reg_9 <= io_host_w_bits_data;
        end
      end
    end
  end
endmodule
module Arbiter( // @[:@178.2]
  output        io_in_0_ready, // @[:@181.4]
  input         io_in_0_valid, // @[:@181.4]
  input  [31:0] io_in_0_bits_addr, // @[:@181.4]
  input  [7:0]  io_in_0_bits_len, // @[:@181.4]
  output        io_in_1_ready, // @[:@181.4]
  input         io_in_1_valid, // @[:@181.4]
  input  [31:0] io_in_1_bits_addr, // @[:@181.4]
  input  [7:0]  io_in_1_bits_len, // @[:@181.4]
  output        io_in_2_ready, // @[:@181.4]
  input         io_in_2_valid, // @[:@181.4]
  input  [31:0] io_in_2_bits_addr, // @[:@181.4]
  input  [7:0]  io_in_2_bits_len, // @[:@181.4]
  output        io_in_3_ready, // @[:@181.4]
  input         io_in_3_valid, // @[:@181.4]
  input  [31:0] io_in_3_bits_addr, // @[:@181.4]
  input  [7:0]  io_in_3_bits_len, // @[:@181.4]
  output        io_in_4_ready, // @[:@181.4]
  input         io_in_4_valid, // @[:@181.4]
  input  [31:0] io_in_4_bits_addr, // @[:@181.4]
  input  [7:0]  io_in_4_bits_len, // @[:@181.4]
  input         io_out_ready, // @[:@181.4]
  output        io_out_valid, // @[:@181.4]
  output [31:0] io_out_bits_addr, // @[:@181.4]
  output [7:0]  io_out_bits_len, // @[:@181.4]
  output [2:0]  io_chosen // @[:@181.4]
);
  wire [2:0] _GEN_0; // @[Arbiter.scala 126:27:@186.4]
  wire [7:0] _GEN_1; // @[Arbiter.scala 126:27:@186.4]
  wire [31:0] _GEN_2; // @[Arbiter.scala 126:27:@186.4]
  wire [2:0] _GEN_3; // @[Arbiter.scala 126:27:@191.4]
  wire [7:0] _GEN_4; // @[Arbiter.scala 126:27:@191.4]
  wire [31:0] _GEN_5; // @[Arbiter.scala 126:27:@191.4]
  wire [2:0] _GEN_6; // @[Arbiter.scala 126:27:@196.4]
  wire [7:0] _GEN_7; // @[Arbiter.scala 126:27:@196.4]
  wire [31:0] _GEN_8; // @[Arbiter.scala 126:27:@196.4]
  wire  _T_114; // @[Arbiter.scala 31:68:@206.4]
  wire  _T_115; // @[Arbiter.scala 31:68:@207.4]
  wire  _T_116; // @[Arbiter.scala 31:68:@208.4]
  wire  _T_118; // @[Arbiter.scala 31:78:@209.4]
  wire  _T_120; // @[Arbiter.scala 31:78:@210.4]
  wire  _T_122; // @[Arbiter.scala 31:78:@211.4]
  wire  _T_124; // @[Arbiter.scala 31:78:@212.4]
  wire  _T_131; // @[Arbiter.scala 135:19:@223.4]
  assign _GEN_0 = io_in_3_valid ? 3'h3 : 3'h4; // @[Arbiter.scala 126:27:@186.4]
  assign _GEN_1 = io_in_3_valid ? io_in_3_bits_len : io_in_4_bits_len; // @[Arbiter.scala 126:27:@186.4]
  assign _GEN_2 = io_in_3_valid ? io_in_3_bits_addr : io_in_4_bits_addr; // @[Arbiter.scala 126:27:@186.4]
  assign _GEN_3 = io_in_2_valid ? 3'h2 : _GEN_0; // @[Arbiter.scala 126:27:@191.4]
  assign _GEN_4 = io_in_2_valid ? io_in_2_bits_len : _GEN_1; // @[Arbiter.scala 126:27:@191.4]
  assign _GEN_5 = io_in_2_valid ? io_in_2_bits_addr : _GEN_2; // @[Arbiter.scala 126:27:@191.4]
  assign _GEN_6 = io_in_1_valid ? 3'h1 : _GEN_3; // @[Arbiter.scala 126:27:@196.4]
  assign _GEN_7 = io_in_1_valid ? io_in_1_bits_len : _GEN_4; // @[Arbiter.scala 126:27:@196.4]
  assign _GEN_8 = io_in_1_valid ? io_in_1_bits_addr : _GEN_5; // @[Arbiter.scala 126:27:@196.4]
  assign _T_114 = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68:@206.4]
  assign _T_115 = _T_114 | io_in_2_valid; // @[Arbiter.scala 31:68:@207.4]
  assign _T_116 = _T_115 | io_in_3_valid; // @[Arbiter.scala 31:68:@208.4]
  assign _T_118 = io_in_0_valid == 1'h0; // @[Arbiter.scala 31:78:@209.4]
  assign _T_120 = _T_114 == 1'h0; // @[Arbiter.scala 31:78:@210.4]
  assign _T_122 = _T_115 == 1'h0; // @[Arbiter.scala 31:78:@211.4]
  assign _T_124 = _T_116 == 1'h0; // @[Arbiter.scala 31:78:@212.4]
  assign _T_131 = _T_124 == 1'h0; // @[Arbiter.scala 135:19:@223.4]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14:@214.4]
  assign io_in_1_ready = _T_118 & io_out_ready; // @[Arbiter.scala 134:14:@216.4]
  assign io_in_2_ready = _T_120 & io_out_ready; // @[Arbiter.scala 134:14:@218.4]
  assign io_in_3_ready = _T_122 & io_out_ready; // @[Arbiter.scala 134:14:@220.4]
  assign io_in_4_ready = _T_124 & io_out_ready; // @[Arbiter.scala 134:14:@222.4]
  assign io_out_valid = _T_131 | io_in_4_valid; // @[Arbiter.scala 135:16:@225.4]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_8; // @[Arbiter.scala 124:15:@185.4 Arbiter.scala 128:19:@189.6 Arbiter.scala 128:19:@194.6 Arbiter.scala 128:19:@199.6 Arbiter.scala 128:19:@204.6]
  assign io_out_bits_len = io_in_0_valid ? io_in_0_bits_len : _GEN_7; // @[Arbiter.scala 124:15:@184.4 Arbiter.scala 128:19:@188.6 Arbiter.scala 128:19:@193.6 Arbiter.scala 128:19:@198.6 Arbiter.scala 128:19:@203.6]
  assign io_chosen = io_in_0_valid ? 3'h0 : _GEN_6; // @[Arbiter.scala 123:13:@183.4 Arbiter.scala 127:17:@187.6 Arbiter.scala 127:17:@192.6 Arbiter.scala 127:17:@197.6 Arbiter.scala 127:17:@202.6]
endmodule
module VME( // @[:@227.2]
  input         clock, // @[:@228.4]
  input         reset, // @[:@229.4]
  input         io_mem_aw_ready, // @[:@230.4]
  output        io_mem_aw_valid, // @[:@230.4]
  output [31:0] io_mem_aw_bits_addr, // @[:@230.4]
  output [7:0]  io_mem_aw_bits_len, // @[:@230.4]
  input         io_mem_w_ready, // @[:@230.4]
  output        io_mem_w_valid, // @[:@230.4]
  output [63:0] io_mem_w_bits_data, // @[:@230.4]
  output        io_mem_w_bits_last, // @[:@230.4]
  output        io_mem_b_ready, // @[:@230.4]
  input         io_mem_b_valid, // @[:@230.4]
  input         io_mem_ar_ready, // @[:@230.4]
  output        io_mem_ar_valid, // @[:@230.4]
  output [31:0] io_mem_ar_bits_addr, // @[:@230.4]
  output [7:0]  io_mem_ar_bits_len, // @[:@230.4]
  output        io_mem_r_ready, // @[:@230.4]
  input         io_mem_r_valid, // @[:@230.4]
  input  [63:0] io_mem_r_bits_data, // @[:@230.4]
  input         io_mem_r_bits_last, // @[:@230.4]
  output        io_vme_rd_0_cmd_ready, // @[:@230.4]
  input         io_vme_rd_0_cmd_valid, // @[:@230.4]
  input  [31:0] io_vme_rd_0_cmd_bits_addr, // @[:@230.4]
  input  [7:0]  io_vme_rd_0_cmd_bits_len, // @[:@230.4]
  input         io_vme_rd_0_data_ready, // @[:@230.4]
  output        io_vme_rd_0_data_valid, // @[:@230.4]
  output [63:0] io_vme_rd_0_data_bits, // @[:@230.4]
  output        io_vme_rd_1_cmd_ready, // @[:@230.4]
  input         io_vme_rd_1_cmd_valid, // @[:@230.4]
  input  [31:0] io_vme_rd_1_cmd_bits_addr, // @[:@230.4]
  input  [7:0]  io_vme_rd_1_cmd_bits_len, // @[:@230.4]
  input         io_vme_rd_1_data_ready, // @[:@230.4]
  output        io_vme_rd_1_data_valid, // @[:@230.4]
  output [63:0] io_vme_rd_1_data_bits, // @[:@230.4]
  output        io_vme_rd_2_cmd_ready, // @[:@230.4]
  input         io_vme_rd_2_cmd_valid, // @[:@230.4]
  input  [31:0] io_vme_rd_2_cmd_bits_addr, // @[:@230.4]
  input  [7:0]  io_vme_rd_2_cmd_bits_len, // @[:@230.4]
  input         io_vme_rd_2_data_ready, // @[:@230.4]
  output        io_vme_rd_2_data_valid, // @[:@230.4]
  output [63:0] io_vme_rd_2_data_bits, // @[:@230.4]
  output        io_vme_rd_3_cmd_ready, // @[:@230.4]
  input         io_vme_rd_3_cmd_valid, // @[:@230.4]
  input  [31:0] io_vme_rd_3_cmd_bits_addr, // @[:@230.4]
  input  [7:0]  io_vme_rd_3_cmd_bits_len, // @[:@230.4]
  input         io_vme_rd_3_data_ready, // @[:@230.4]
  output        io_vme_rd_3_data_valid, // @[:@230.4]
  output [63:0] io_vme_rd_3_data_bits, // @[:@230.4]
  output        io_vme_rd_4_cmd_ready, // @[:@230.4]
  input         io_vme_rd_4_cmd_valid, // @[:@230.4]
  input  [31:0] io_vme_rd_4_cmd_bits_addr, // @[:@230.4]
  input  [7:0]  io_vme_rd_4_cmd_bits_len, // @[:@230.4]
  input         io_vme_rd_4_data_ready, // @[:@230.4]
  output        io_vme_rd_4_data_valid, // @[:@230.4]
  output [63:0] io_vme_rd_4_data_bits, // @[:@230.4]
  output        io_vme_wr_0_cmd_ready, // @[:@230.4]
  input         io_vme_wr_0_cmd_valid, // @[:@230.4]
  input  [31:0] io_vme_wr_0_cmd_bits_addr, // @[:@230.4]
  input  [7:0]  io_vme_wr_0_cmd_bits_len, // @[:@230.4]
  output        io_vme_wr_0_data_ready, // @[:@230.4]
  input         io_vme_wr_0_data_valid, // @[:@230.4]
  input  [63:0] io_vme_wr_0_data_bits, // @[:@230.4]
  output        io_vme_wr_0_ack // @[:@230.4]
);
  wire  rd_arb_io_in_0_ready; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_in_0_valid; // @[VME.scala 146:22:@232.4]
  wire [31:0] rd_arb_io_in_0_bits_addr; // @[VME.scala 146:22:@232.4]
  wire [7:0] rd_arb_io_in_0_bits_len; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_in_1_ready; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_in_1_valid; // @[VME.scala 146:22:@232.4]
  wire [31:0] rd_arb_io_in_1_bits_addr; // @[VME.scala 146:22:@232.4]
  wire [7:0] rd_arb_io_in_1_bits_len; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_in_2_ready; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_in_2_valid; // @[VME.scala 146:22:@232.4]
  wire [31:0] rd_arb_io_in_2_bits_addr; // @[VME.scala 146:22:@232.4]
  wire [7:0] rd_arb_io_in_2_bits_len; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_in_3_ready; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_in_3_valid; // @[VME.scala 146:22:@232.4]
  wire [31:0] rd_arb_io_in_3_bits_addr; // @[VME.scala 146:22:@232.4]
  wire [7:0] rd_arb_io_in_3_bits_len; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_in_4_ready; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_in_4_valid; // @[VME.scala 146:22:@232.4]
  wire [31:0] rd_arb_io_in_4_bits_addr; // @[VME.scala 146:22:@232.4]
  wire [7:0] rd_arb_io_in_4_bits_len; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_out_ready; // @[VME.scala 146:22:@232.4]
  wire  rd_arb_io_out_valid; // @[VME.scala 146:22:@232.4]
  wire [31:0] rd_arb_io_out_bits_addr; // @[VME.scala 146:22:@232.4]
  wire [7:0] rd_arb_io_out_bits_len; // @[VME.scala 146:22:@232.4]
  wire [2:0] rd_arb_io_chosen; // @[VME.scala 146:22:@232.4]
  wire  _T_260; // @[Decoupled.scala 37:37:@235.4]
  reg [2:0] rd_arb_chosen; // @[Reg.scala 11:16:@236.4]
  reg [31:0] _RAND_0;
  reg [1:0] rstate; // @[VME.scala 152:23:@260.4]
  reg [31:0] _RAND_1;
  wire  _T_263; // @[Conditional.scala 37:30:@261.4]
  wire [1:0] _GEN_1; // @[VME.scala 156:33:@263.6]
  wire  _T_264; // @[Conditional.scala 37:30:@268.6]
  wire [1:0] _GEN_2; // @[VME.scala 161:29:@270.8]
  wire  _T_265; // @[Conditional.scala 37:30:@275.8]
  wire  _T_266; // @[Decoupled.scala 37:37:@277.10]
  wire  _T_267; // @[VME.scala 166:28:@278.10]
  wire [1:0] _GEN_3; // @[VME.scala 166:51:@279.10]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@276.8]
  wire [1:0] _GEN_5; // @[Conditional.scala 39:67:@269.6]
  wire [1:0] _GEN_6; // @[Conditional.scala 40:58:@262.4]
  reg [1:0] wstate; // @[VME.scala 173:23:@283.4]
  reg [31:0] _RAND_2;
  reg [7:0] wr_cnt; // @[VME.scala 176:23:@284.4]
  reg [31:0] _RAND_3;
  wire  _T_271; // @[VME.scala 178:15:@285.4]
  wire  _T_273; // @[Decoupled.scala 37:37:@290.6]
  wire [8:0] _T_275; // @[VME.scala 181:22:@292.8]
  wire [7:0] _T_276; // @[VME.scala 181:22:@293.8]
  wire [7:0] _GEN_7; // @[VME.scala 180:31:@291.6]
  wire [7:0] _GEN_8; // @[VME.scala 178:31:@286.4]
  wire  _T_277; // @[Conditional.scala 37:30:@296.4]
  wire [1:0] _GEN_9; // @[VME.scala 186:36:@298.6]
  wire  _T_278; // @[Conditional.scala 37:30:@303.6]
  wire [1:0] _GEN_10; // @[VME.scala 191:29:@305.8]
  wire  _T_279; // @[Conditional.scala 37:30:@310.8]
  wire  _T_280; // @[VME.scala 200:18:@312.10]
  wire  _T_281; // @[VME.scala 200:46:@313.10]
  wire  _T_282; // @[VME.scala 200:36:@314.10]
  wire [1:0] _GEN_11; // @[VME.scala 200:77:@315.10]
  wire  _T_283; // @[Conditional.scala 37:30:@320.10]
  wire [1:0] _GEN_12; // @[VME.scala 205:28:@322.12]
  wire [1:0] _GEN_13; // @[Conditional.scala 39:67:@321.10]
  wire [1:0] _GEN_14; // @[Conditional.scala 39:67:@311.8]
  wire [1:0] _GEN_15; // @[Conditional.scala 39:67:@304.6]
  wire [1:0] _GEN_16; // @[Conditional.scala 40:58:@297.4]
  reg [7:0] rd_len; // @[VME.scala 213:23:@326.4]
  reg [31:0] _RAND_4;
  reg [7:0] wr_len; // @[VME.scala 214:23:@327.4]
  reg [31:0] _RAND_5;
  reg [31:0] rd_addr; // @[VME.scala 215:24:@328.4]
  reg [31:0] _RAND_6;
  reg [31:0] wr_addr; // @[VME.scala 216:24:@329.4]
  reg [31:0] _RAND_7;
  wire [7:0] _GEN_17; // @[VME.scala 218:30:@331.4]
  wire [31:0] _GEN_18; // @[VME.scala 218:30:@331.4]
  wire  _T_293; // @[Decoupled.scala 37:37:@335.4]
  wire [7:0] _GEN_19; // @[VME.scala 223:33:@336.4]
  wire [31:0] _GEN_20; // @[VME.scala 223:33:@336.4]
  wire  _T_296; // @[VME.scala 233:46:@342.4]
  wire  _T_299; // @[VME.scala 233:46:@346.4]
  wire  _T_302; // @[VME.scala 233:46:@350.4]
  wire  _T_305; // @[VME.scala 233:46:@354.4]
  wire  _T_308; // @[VME.scala 233:46:@358.4]
  wire  _T_312; // @[VME.scala 239:37:@366.4]
  wire  _T_320; // @[VME.scala 256:28:@385.4]
  wire  _GEN_32; // @[VME.scala 256:42:@386.4]
  wire  _GEN_39; // @[VME.scala 256:42:@386.4]
  wire  _GEN_46; // @[VME.scala 256:42:@386.4]
  wire  _GEN_53; // @[VME.scala 256:42:@386.4]
  Arbiter rd_arb ( // @[VME.scala 146:22:@232.4]
    .io_in_0_ready(rd_arb_io_in_0_ready),
    .io_in_0_valid(rd_arb_io_in_0_valid),
    .io_in_0_bits_addr(rd_arb_io_in_0_bits_addr),
    .io_in_0_bits_len(rd_arb_io_in_0_bits_len),
    .io_in_1_ready(rd_arb_io_in_1_ready),
    .io_in_1_valid(rd_arb_io_in_1_valid),
    .io_in_1_bits_addr(rd_arb_io_in_1_bits_addr),
    .io_in_1_bits_len(rd_arb_io_in_1_bits_len),
    .io_in_2_ready(rd_arb_io_in_2_ready),
    .io_in_2_valid(rd_arb_io_in_2_valid),
    .io_in_2_bits_addr(rd_arb_io_in_2_bits_addr),
    .io_in_2_bits_len(rd_arb_io_in_2_bits_len),
    .io_in_3_ready(rd_arb_io_in_3_ready),
    .io_in_3_valid(rd_arb_io_in_3_valid),
    .io_in_3_bits_addr(rd_arb_io_in_3_bits_addr),
    .io_in_3_bits_len(rd_arb_io_in_3_bits_len),
    .io_in_4_ready(rd_arb_io_in_4_ready),
    .io_in_4_valid(rd_arb_io_in_4_valid),
    .io_in_4_bits_addr(rd_arb_io_in_4_bits_addr),
    .io_in_4_bits_len(rd_arb_io_in_4_bits_len),
    .io_out_ready(rd_arb_io_out_ready),
    .io_out_valid(rd_arb_io_out_valid),
    .io_out_bits_addr(rd_arb_io_out_bits_addr),
    .io_out_bits_len(rd_arb_io_out_bits_len),
    .io_chosen(rd_arb_io_chosen)
  );
  assign _T_260 = rd_arb_io_out_ready & rd_arb_io_out_valid; // @[Decoupled.scala 37:37:@235.4]
  assign _T_263 = 2'h0 == rstate; // @[Conditional.scala 37:30:@261.4]
  assign _GEN_1 = rd_arb_io_out_valid ? 2'h1 : rstate; // @[VME.scala 156:33:@263.6]
  assign _T_264 = 2'h1 == rstate; // @[Conditional.scala 37:30:@268.6]
  assign _GEN_2 = io_mem_ar_ready ? 2'h2 : rstate; // @[VME.scala 161:29:@270.8]
  assign _T_265 = 2'h2 == rstate; // @[Conditional.scala 37:30:@275.8]
  assign _T_266 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 37:37:@277.10]
  assign _T_267 = _T_266 & io_mem_r_bits_last; // @[VME.scala 166:28:@278.10]
  assign _GEN_3 = _T_267 ? 2'h0 : rstate; // @[VME.scala 166:51:@279.10]
  assign _GEN_4 = _T_265 ? _GEN_3 : rstate; // @[Conditional.scala 39:67:@276.8]
  assign _GEN_5 = _T_264 ? _GEN_2 : _GEN_4; // @[Conditional.scala 39:67:@269.6]
  assign _GEN_6 = _T_263 ? _GEN_1 : _GEN_5; // @[Conditional.scala 40:58:@262.4]
  assign _T_271 = wstate == 2'h0; // @[VME.scala 178:15:@285.4]
  assign _T_273 = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 37:37:@290.6]
  assign _T_275 = wr_cnt + 8'h1; // @[VME.scala 181:22:@292.8]
  assign _T_276 = wr_cnt + 8'h1; // @[VME.scala 181:22:@293.8]
  assign _GEN_7 = _T_273 ? _T_276 : wr_cnt; // @[VME.scala 180:31:@291.6]
  assign _GEN_8 = _T_271 ? 8'h0 : _GEN_7; // @[VME.scala 178:31:@286.4]
  assign _T_277 = 2'h0 == wstate; // @[Conditional.scala 37:30:@296.4]
  assign _GEN_9 = io_vme_wr_0_cmd_valid ? 2'h1 : wstate; // @[VME.scala 186:36:@298.6]
  assign _T_278 = 2'h1 == wstate; // @[Conditional.scala 37:30:@303.6]
  assign _GEN_10 = io_mem_aw_ready ? 2'h2 : wstate; // @[VME.scala 191:29:@305.8]
  assign _T_279 = 2'h2 == wstate; // @[Conditional.scala 37:30:@310.8]
  assign _T_280 = io_vme_wr_0_data_valid & io_mem_w_ready; // @[VME.scala 200:18:@312.10]
  assign _T_281 = wr_cnt == io_vme_wr_0_cmd_bits_len; // @[VME.scala 200:46:@313.10]
  assign _T_282 = _T_280 & _T_281; // @[VME.scala 200:36:@314.10]
  assign _GEN_11 = _T_282 ? 2'h3 : wstate; // @[VME.scala 200:77:@315.10]
  assign _T_283 = 2'h3 == wstate; // @[Conditional.scala 37:30:@320.10]
  assign _GEN_12 = io_mem_b_valid ? 2'h0 : wstate; // @[VME.scala 205:28:@322.12]
  assign _GEN_13 = _T_283 ? _GEN_12 : wstate; // @[Conditional.scala 39:67:@321.10]
  assign _GEN_14 = _T_279 ? _GEN_11 : _GEN_13; // @[Conditional.scala 39:67:@311.8]
  assign _GEN_15 = _T_278 ? _GEN_10 : _GEN_14; // @[Conditional.scala 39:67:@304.6]
  assign _GEN_16 = _T_277 ? _GEN_9 : _GEN_15; // @[Conditional.scala 40:58:@297.4]
  assign _GEN_17 = _T_260 ? rd_arb_io_out_bits_len : rd_len; // @[VME.scala 218:30:@331.4]
  assign _GEN_18 = _T_260 ? rd_arb_io_out_bits_addr : rd_addr; // @[VME.scala 218:30:@331.4]
  assign _T_293 = io_vme_wr_0_cmd_ready & io_vme_wr_0_cmd_valid; // @[Decoupled.scala 37:37:@335.4]
  assign _GEN_19 = _T_293 ? io_vme_wr_0_cmd_bits_len : wr_len; // @[VME.scala 223:33:@336.4]
  assign _GEN_20 = _T_293 ? io_vme_wr_0_cmd_bits_addr : wr_addr; // @[VME.scala 223:33:@336.4]
  assign _T_296 = rd_arb_chosen == 3'h0; // @[VME.scala 233:46:@342.4]
  assign _T_299 = rd_arb_chosen == 3'h1; // @[VME.scala 233:46:@346.4]
  assign _T_302 = rd_arb_chosen == 3'h2; // @[VME.scala 233:46:@350.4]
  assign _T_305 = rd_arb_chosen == 3'h3; // @[VME.scala 233:46:@354.4]
  assign _T_308 = rd_arb_chosen == 3'h4; // @[VME.scala 233:46:@358.4]
  assign _T_312 = wstate == 2'h2; // @[VME.scala 239:37:@366.4]
  assign _T_320 = rstate == 2'h2; // @[VME.scala 256:28:@385.4]
  assign _GEN_32 = 3'h1 == rd_arb_chosen ? io_vme_rd_1_data_ready : io_vme_rd_0_data_ready; // @[VME.scala 256:42:@386.4]
  assign _GEN_39 = 3'h2 == rd_arb_chosen ? io_vme_rd_2_data_ready : _GEN_32; // @[VME.scala 256:42:@386.4]
  assign _GEN_46 = 3'h3 == rd_arb_chosen ? io_vme_rd_3_data_ready : _GEN_39; // @[VME.scala 256:42:@386.4]
  assign _GEN_53 = 3'h4 == rd_arb_chosen ? io_vme_rd_4_data_ready : _GEN_46; // @[VME.scala 256:42:@386.4]
  assign io_mem_aw_valid = wstate == 2'h1; // @[VME.scala 242:19:@370.4]
  assign io_mem_aw_bits_addr = wr_addr; // @[VME.scala 243:23:@371.4]
  assign io_mem_aw_bits_len = wr_len; // @[VME.scala 244:22:@372.4]
  assign io_mem_w_valid = _T_312 & io_vme_wr_0_data_valid; // @[VME.scala 246:18:@375.4]
  assign io_mem_w_bits_data = io_vme_wr_0_data_bits; // @[VME.scala 247:22:@376.4]
  assign io_mem_w_bits_last = wr_cnt == io_vme_wr_0_cmd_bits_len; // @[VME.scala 248:22:@378.4]
  assign io_mem_b_ready = wstate == 2'h3; // @[VME.scala 250:18:@380.4]
  assign io_mem_ar_valid = rstate == 2'h1; // @[VME.scala 252:19:@382.4]
  assign io_mem_ar_bits_addr = rd_addr; // @[VME.scala 253:23:@383.4]
  assign io_mem_ar_bits_len = rd_len; // @[VME.scala 254:22:@384.4]
  assign io_mem_r_ready = _T_320 & _GEN_53; // @[VME.scala 256:18:@387.4]
  assign io_vme_rd_0_cmd_ready = rd_arb_io_in_0_ready; // @[VME.scala 149:53:@243.4]
  assign io_vme_rd_0_data_valid = _T_296 & io_mem_r_valid; // @[VME.scala 233:29:@344.4]
  assign io_vme_rd_0_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@345.4]
  assign io_vme_rd_1_cmd_ready = rd_arb_io_in_1_ready; // @[VME.scala 149:53:@247.4]
  assign io_vme_rd_1_data_valid = _T_299 & io_mem_r_valid; // @[VME.scala 233:29:@348.4]
  assign io_vme_rd_1_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@349.4]
  assign io_vme_rd_2_cmd_ready = rd_arb_io_in_2_ready; // @[VME.scala 149:53:@251.4]
  assign io_vme_rd_2_data_valid = _T_302 & io_mem_r_valid; // @[VME.scala 233:29:@352.4]
  assign io_vme_rd_2_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@353.4]
  assign io_vme_rd_3_cmd_ready = rd_arb_io_in_3_ready; // @[VME.scala 149:53:@255.4]
  assign io_vme_rd_3_data_valid = _T_305 & io_mem_r_valid; // @[VME.scala 233:29:@356.4]
  assign io_vme_rd_3_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@357.4]
  assign io_vme_rd_4_cmd_ready = rd_arb_io_in_4_ready; // @[VME.scala 149:53:@259.4]
  assign io_vme_rd_4_data_valid = _T_308 & io_mem_r_valid; // @[VME.scala 233:29:@360.4]
  assign io_vme_rd_4_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@361.4]
  assign io_vme_wr_0_cmd_ready = wstate == 2'h0; // @[VME.scala 237:26:@363.4]
  assign io_vme_wr_0_data_ready = _T_312 & io_mem_w_ready; // @[VME.scala 239:27:@368.4]
  assign io_vme_wr_0_ack = io_mem_b_ready & io_mem_b_valid; // @[VME.scala 238:20:@365.4]
  assign rd_arb_io_in_0_valid = io_vme_rd_0_cmd_valid; // @[VME.scala 149:53:@242.4]
  assign rd_arb_io_in_0_bits_addr = io_vme_rd_0_cmd_bits_addr; // @[VME.scala 149:53:@241.4]
  assign rd_arb_io_in_0_bits_len = io_vme_rd_0_cmd_bits_len; // @[VME.scala 149:53:@240.4]
  assign rd_arb_io_in_1_valid = io_vme_rd_1_cmd_valid; // @[VME.scala 149:53:@246.4]
  assign rd_arb_io_in_1_bits_addr = io_vme_rd_1_cmd_bits_addr; // @[VME.scala 149:53:@245.4]
  assign rd_arb_io_in_1_bits_len = io_vme_rd_1_cmd_bits_len; // @[VME.scala 149:53:@244.4]
  assign rd_arb_io_in_2_valid = io_vme_rd_2_cmd_valid; // @[VME.scala 149:53:@250.4]
  assign rd_arb_io_in_2_bits_addr = io_vme_rd_2_cmd_bits_addr; // @[VME.scala 149:53:@249.4]
  assign rd_arb_io_in_2_bits_len = io_vme_rd_2_cmd_bits_len; // @[VME.scala 149:53:@248.4]
  assign rd_arb_io_in_3_valid = io_vme_rd_3_cmd_valid; // @[VME.scala 149:53:@254.4]
  assign rd_arb_io_in_3_bits_addr = io_vme_rd_3_cmd_bits_addr; // @[VME.scala 149:53:@253.4]
  assign rd_arb_io_in_3_bits_len = io_vme_rd_3_cmd_bits_len; // @[VME.scala 149:53:@252.4]
  assign rd_arb_io_in_4_valid = io_vme_rd_4_cmd_valid; // @[VME.scala 149:53:@258.4]
  assign rd_arb_io_in_4_bits_addr = io_vme_rd_4_cmd_bits_addr; // @[VME.scala 149:53:@257.4]
  assign rd_arb_io_in_4_bits_len = io_vme_rd_4_cmd_bits_len; // @[VME.scala 149:53:@256.4]
  assign rd_arb_io_out_ready = rstate == 2'h0; // @[VME.scala 229:23:@341.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_arb_chosen = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rstate = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  wstate = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  wr_cnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_len = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  wr_len = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  wr_addr = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_260) begin
      rd_arb_chosen <= rd_arb_io_chosen;
    end
    if (reset) begin
      rstate <= 2'h0;
    end else begin
      if (_T_263) begin
        if (rd_arb_io_out_valid) begin
          rstate <= 2'h1;
        end
      end else begin
        if (_T_264) begin
          if (io_mem_ar_ready) begin
            rstate <= 2'h2;
          end
        end else begin
          if (_T_265) begin
            if (_T_267) begin
              rstate <= 2'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      wstate <= 2'h0;
    end else begin
      if (_T_277) begin
        if (io_vme_wr_0_cmd_valid) begin
          wstate <= 2'h1;
        end
      end else begin
        if (_T_278) begin
          if (io_mem_aw_ready) begin
            wstate <= 2'h2;
          end
        end else begin
          if (_T_279) begin
            if (_T_282) begin
              wstate <= 2'h3;
            end
          end else begin
            if (_T_283) begin
              if (io_mem_b_valid) begin
                wstate <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      wr_cnt <= 8'h0;
    end else begin
      if (_T_271) begin
        wr_cnt <= 8'h0;
      end else begin
        if (_T_273) begin
          wr_cnt <= _T_276;
        end
      end
    end
    if (reset) begin
      rd_len <= 8'h0;
    end else begin
      if (_T_260) begin
        rd_len <= rd_arb_io_out_bits_len;
      end
    end
    if (reset) begin
      wr_len <= 8'h0;
    end else begin
      if (_T_293) begin
        wr_len <= io_vme_wr_0_cmd_bits_len;
      end
    end
    if (reset) begin
      rd_addr <= 32'h0;
    end else begin
      if (_T_260) begin
        rd_addr <= rd_arb_io_out_bits_addr;
      end
    end
    if (reset) begin
      wr_addr <= 32'h0;
    end else begin
      if (_T_293) begin
        wr_addr <= io_vme_wr_0_cmd_bits_addr;
      end
    end
  end
endmodule
module Queue( // @[:@411.2]
  input          clock, // @[:@412.4]
  input          reset, // @[:@413.4]
  output         io_enq_ready, // @[:@414.4]
  input          io_enq_valid, // @[:@414.4]
  input  [127:0] io_enq_bits, // @[:@414.4]
  input          io_deq_ready, // @[:@414.4]
  output         io_deq_valid, // @[:@414.4]
  output [127:0] io_deq_bits, // @[:@414.4]
  output [7:0]   io_count // @[:@414.4]
);
  reg [127:0] _T_35 [0:127]; // @[Decoupled.scala 215:24:@416.4]
  reg [127:0] _RAND_0;
  wire [127:0] _T_35__T_68_data; // @[Decoupled.scala 215:24:@416.4]
  wire [6:0] _T_35__T_68_addr; // @[Decoupled.scala 215:24:@416.4]
  wire [127:0] _T_35__T_54_data; // @[Decoupled.scala 215:24:@416.4]
  wire [6:0] _T_35__T_54_addr; // @[Decoupled.scala 215:24:@416.4]
  wire  _T_35__T_54_mask; // @[Decoupled.scala 215:24:@416.4]
  wire  _T_35__T_54_en; // @[Decoupled.scala 215:24:@416.4]
  reg [6:0] value; // @[Counter.scala 26:33:@417.4]
  reg [31:0] _RAND_1;
  reg [6:0] value_1; // @[Counter.scala 26:33:@418.4]
  reg [31:0] _RAND_2;
  reg  _T_42; // @[Decoupled.scala 218:35:@419.4]
  reg [31:0] _RAND_3;
  wire  _T_43; // @[Decoupled.scala 220:41:@420.4]
  wire  _T_45; // @[Decoupled.scala 221:36:@421.4]
  wire  _T_46; // @[Decoupled.scala 221:33:@422.4]
  wire  _T_47; // @[Decoupled.scala 222:32:@423.4]
  wire  _T_48; // @[Decoupled.scala 37:37:@424.4]
  wire  _T_51; // @[Decoupled.scala 37:37:@427.4]
  wire [7:0] _T_57; // @[Counter.scala 35:22:@434.6]
  wire [6:0] _T_58; // @[Counter.scala 35:22:@435.6]
  wire [6:0] _GEN_5; // @[Decoupled.scala 226:17:@430.4]
  wire [7:0] _T_61; // @[Counter.scala 35:22:@440.6]
  wire [6:0] _T_62; // @[Counter.scala 35:22:@441.6]
  wire [6:0] _GEN_6; // @[Decoupled.scala 230:17:@438.4]
  wire  _T_63; // @[Decoupled.scala 233:16:@444.4]
  wire  _GEN_7; // @[Decoupled.scala 233:28:@445.4]
  wire [7:0] _T_69; // @[Decoupled.scala 254:40:@454.4]
  wire [7:0] _T_70; // @[Decoupled.scala 254:40:@455.4]
  wire [6:0] _T_71; // @[Decoupled.scala 254:40:@456.4]
  wire  _T_72; // @[Decoupled.scala 256:32:@457.4]
  wire [7:0] _T_75; // @[Decoupled.scala 256:20:@458.4]
  wire [7:0] _GEN_14; // @[Decoupled.scala 256:62:@459.4]
  assign _T_35__T_68_addr = value_1;
  assign _T_35__T_68_data = _T_35[_T_35__T_68_addr]; // @[Decoupled.scala 215:24:@416.4]
  assign _T_35__T_54_data = io_enq_bits;
  assign _T_35__T_54_addr = value;
  assign _T_35__T_54_mask = 1'h1;
  assign _T_35__T_54_en = io_enq_ready & io_enq_valid;
  assign _T_43 = value == value_1; // @[Decoupled.scala 220:41:@420.4]
  assign _T_45 = _T_42 == 1'h0; // @[Decoupled.scala 221:36:@421.4]
  assign _T_46 = _T_43 & _T_45; // @[Decoupled.scala 221:33:@422.4]
  assign _T_47 = _T_43 & _T_42; // @[Decoupled.scala 222:32:@423.4]
  assign _T_48 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:@424.4]
  assign _T_51 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:@427.4]
  assign _T_57 = value + 7'h1; // @[Counter.scala 35:22:@434.6]
  assign _T_58 = value + 7'h1; // @[Counter.scala 35:22:@435.6]
  assign _GEN_5 = _T_48 ? _T_58 : value; // @[Decoupled.scala 226:17:@430.4]
  assign _T_61 = value_1 + 7'h1; // @[Counter.scala 35:22:@440.6]
  assign _T_62 = value_1 + 7'h1; // @[Counter.scala 35:22:@441.6]
  assign _GEN_6 = _T_51 ? _T_62 : value_1; // @[Decoupled.scala 230:17:@438.4]
  assign _T_63 = _T_48 != _T_51; // @[Decoupled.scala 233:16:@444.4]
  assign _GEN_7 = _T_63 ? _T_48 : _T_42; // @[Decoupled.scala 233:28:@445.4]
  assign _T_69 = value - value_1; // @[Decoupled.scala 254:40:@454.4]
  assign _T_70 = $unsigned(_T_69); // @[Decoupled.scala 254:40:@455.4]
  assign _T_71 = _T_70[6:0]; // @[Decoupled.scala 254:40:@456.4]
  assign _T_72 = _T_42 & _T_43; // @[Decoupled.scala 256:32:@457.4]
  assign _T_75 = _T_72 ? 8'h80 : 8'h0; // @[Decoupled.scala 256:20:@458.4]
  assign _GEN_14 = {{1'd0}, _T_71}; // @[Decoupled.scala 256:62:@459.4]
  assign io_enq_ready = _T_47 == 1'h0; // @[Decoupled.scala 238:16:@451.4]
  assign io_deq_valid = _T_46 == 1'h0; // @[Decoupled.scala 237:16:@449.4]
  assign io_deq_bits = _T_35__T_68_data; // @[Decoupled.scala 239:15:@453.4]
  assign io_count = _T_75 | _GEN_14; // @[Decoupled.scala 256:14:@460.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T_35[initvar] = _RAND_0[127:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_42 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35__T_54_en & _T_35__T_54_mask) begin
      _T_35[_T_35__T_54_addr] <= _T_35__T_54_data; // @[Decoupled.scala 215:24:@416.4]
    end
    if (reset) begin
      value <= 7'h0;
    end else begin
      if (_T_48) begin
        value <= _T_58;
      end
    end
    if (reset) begin
      value_1 <= 7'h0;
    end else begin
      if (_T_51) begin
        value_1 <= _T_62;
      end
    end
    if (reset) begin
      _T_42 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_42 <= _T_48;
      end
    end
  end
endmodule
module FetchDecode( // @[:@462.2]
  input  [127:0] io_inst, // @[:@465.4]
  output         io_isLoad, // @[:@465.4]
  output         io_isCompute, // @[:@465.4]
  output         io_isStore // @[:@465.4]
);
  wire [127:0] _T_15; // @[Lookup.scala 9:38:@467.4]
  wire  _T_16; // @[Lookup.scala 9:38:@468.4]
  wire  _T_20; // @[Lookup.scala 9:38:@470.4]
  wire  _T_24; // @[Lookup.scala 9:38:@472.4]
  wire  _T_28; // @[Lookup.scala 9:38:@474.4]
  wire [127:0] _T_31; // @[Lookup.scala 9:38:@475.4]
  wire  _T_32; // @[Lookup.scala 9:38:@476.4]
  wire  _T_36; // @[Lookup.scala 9:38:@478.4]
  wire  _T_40; // @[Lookup.scala 9:38:@480.4]
  wire [127:0] _T_43; // @[Lookup.scala 9:38:@481.4]
  wire  _T_44; // @[Lookup.scala 9:38:@482.4]
  wire  _T_48; // @[Lookup.scala 9:38:@484.4]
  wire  _T_52; // @[Lookup.scala 9:38:@486.4]
  wire  _T_56; // @[Lookup.scala 9:38:@488.4]
  wire  _T_58; // @[Lookup.scala 11:37:@490.4]
  wire  _T_59; // @[Lookup.scala 11:37:@491.4]
  wire  _T_60; // @[Lookup.scala 11:37:@492.4]
  wire  _T_61; // @[Lookup.scala 11:37:@493.4]
  wire  _T_62; // @[Lookup.scala 11:37:@494.4]
  wire  _T_63; // @[Lookup.scala 11:37:@495.4]
  wire  _T_64; // @[Lookup.scala 11:37:@496.4]
  wire  _T_65; // @[Lookup.scala 11:37:@497.4]
  wire  _T_66; // @[Lookup.scala 11:37:@498.4]
  wire  cs_val_inst; // @[Lookup.scala 11:37:@499.4]
  wire [2:0] _T_67; // @[Lookup.scala 11:37:@500.4]
  wire [2:0] _T_68; // @[Lookup.scala 11:37:@501.4]
  wire [2:0] _T_69; // @[Lookup.scala 11:37:@502.4]
  wire [2:0] _T_70; // @[Lookup.scala 11:37:@503.4]
  wire [2:0] _T_71; // @[Lookup.scala 11:37:@504.4]
  wire [2:0] _T_72; // @[Lookup.scala 11:37:@505.4]
  wire [2:0] _T_73; // @[Lookup.scala 11:37:@506.4]
  wire [2:0] _T_74; // @[Lookup.scala 11:37:@507.4]
  wire [2:0] _T_75; // @[Lookup.scala 11:37:@508.4]
  wire [2:0] _T_76; // @[Lookup.scala 11:37:@509.4]
  wire [2:0] cs_op_type; // @[Lookup.scala 11:37:@510.4]
  wire  _T_77; // @[Decode.scala 156:41:@511.4]
  wire  _T_79; // @[Decode.scala 157:44:@514.4]
  wire  _T_81; // @[Decode.scala 158:42:@517.4]
  assign _T_15 = io_inst & 128'h187; // @[Lookup.scala 9:38:@467.4]
  assign _T_16 = 128'h0 == _T_15; // @[Lookup.scala 9:38:@468.4]
  assign _T_20 = 128'h80 == _T_15; // @[Lookup.scala 9:38:@470.4]
  assign _T_24 = 128'h100 == _T_15; // @[Lookup.scala 9:38:@472.4]
  assign _T_28 = 128'h180 == _T_15; // @[Lookup.scala 9:38:@474.4]
  assign _T_31 = io_inst & 128'h7; // @[Lookup.scala 9:38:@475.4]
  assign _T_32 = 128'h1 == _T_31; // @[Lookup.scala 9:38:@476.4]
  assign _T_36 = 128'h2 == _T_31; // @[Lookup.scala 9:38:@478.4]
  assign _T_40 = 128'h3 == _T_31; // @[Lookup.scala 9:38:@480.4]
  assign _T_43 = io_inst & 128'h3000000000000000000000000007; // @[Lookup.scala 9:38:@481.4]
  assign _T_44 = 128'h4 == _T_43; // @[Lookup.scala 9:38:@482.4]
  assign _T_48 = 128'h1000000000000000000000000004 == _T_43; // @[Lookup.scala 9:38:@484.4]
  assign _T_52 = 128'h2000000000000000000000000004 == _T_43; // @[Lookup.scala 9:38:@486.4]
  assign _T_56 = 128'h3000000000000000000000000004 == _T_43; // @[Lookup.scala 9:38:@488.4]
  assign _T_58 = _T_52 ? 1'h1 : _T_56; // @[Lookup.scala 11:37:@490.4]
  assign _T_59 = _T_48 ? 1'h1 : _T_58; // @[Lookup.scala 11:37:@491.4]
  assign _T_60 = _T_44 ? 1'h1 : _T_59; // @[Lookup.scala 11:37:@492.4]
  assign _T_61 = _T_40 ? 1'h1 : _T_60; // @[Lookup.scala 11:37:@493.4]
  assign _T_62 = _T_36 ? 1'h1 : _T_61; // @[Lookup.scala 11:37:@494.4]
  assign _T_63 = _T_32 ? 1'h1 : _T_62; // @[Lookup.scala 11:37:@495.4]
  assign _T_64 = _T_28 ? 1'h1 : _T_63; // @[Lookup.scala 11:37:@496.4]
  assign _T_65 = _T_24 ? 1'h1 : _T_64; // @[Lookup.scala 11:37:@497.4]
  assign _T_66 = _T_20 ? 1'h1 : _T_65; // @[Lookup.scala 11:37:@498.4]
  assign cs_val_inst = _T_16 ? 1'h1 : _T_66; // @[Lookup.scala 11:37:@499.4]
  assign _T_67 = _T_56 ? 3'h2 : 3'h5; // @[Lookup.scala 11:37:@500.4]
  assign _T_68 = _T_52 ? 3'h2 : _T_67; // @[Lookup.scala 11:37:@501.4]
  assign _T_69 = _T_48 ? 3'h2 : _T_68; // @[Lookup.scala 11:37:@502.4]
  assign _T_70 = _T_44 ? 3'h2 : _T_69; // @[Lookup.scala 11:37:@503.4]
  assign _T_71 = _T_40 ? 3'h2 : _T_70; // @[Lookup.scala 11:37:@504.4]
  assign _T_72 = _T_36 ? 3'h2 : _T_71; // @[Lookup.scala 11:37:@505.4]
  assign _T_73 = _T_32 ? 3'h1 : _T_72; // @[Lookup.scala 11:37:@506.4]
  assign _T_74 = _T_28 ? 3'h2 : _T_73; // @[Lookup.scala 11:37:@507.4]
  assign _T_75 = _T_24 ? 3'h0 : _T_74; // @[Lookup.scala 11:37:@508.4]
  assign _T_76 = _T_20 ? 3'h0 : _T_75; // @[Lookup.scala 11:37:@509.4]
  assign cs_op_type = _T_16 ? 3'h2 : _T_76; // @[Lookup.scala 11:37:@510.4]
  assign _T_77 = cs_op_type == 3'h0; // @[Decode.scala 156:41:@511.4]
  assign _T_79 = cs_op_type == 3'h2; // @[Decode.scala 157:44:@514.4]
  assign _T_81 = cs_op_type == 3'h1; // @[Decode.scala 158:42:@517.4]
  assign io_isLoad = cs_val_inst & _T_77; // @[Decode.scala 156:13:@513.4]
  assign io_isCompute = cs_val_inst & _T_79; // @[Decode.scala 157:16:@516.4]
  assign io_isStore = cs_val_inst & _T_81; // @[Decode.scala 158:14:@519.4]
endmodule
module Fetch( // @[:@521.2]
  input          clock, // @[:@522.4]
  input          reset, // @[:@523.4]
  input          io_launch, // @[:@524.4]
  input  [31:0]  io_ins_baddr, // @[:@524.4]
  input  [31:0]  io_ins_count, // @[:@524.4]
  input          io_vme_rd_cmd_ready, // @[:@524.4]
  output         io_vme_rd_cmd_valid, // @[:@524.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@524.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@524.4]
  output         io_vme_rd_data_ready, // @[:@524.4]
  input          io_vme_rd_data_valid, // @[:@524.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@524.4]
  input          io_inst_ld_ready, // @[:@524.4]
  output         io_inst_ld_valid, // @[:@524.4]
  output [127:0] io_inst_ld_bits, // @[:@524.4]
  input          io_inst_co_ready, // @[:@524.4]
  output         io_inst_co_valid, // @[:@524.4]
  output [127:0] io_inst_co_bits, // @[:@524.4]
  input          io_inst_st_ready, // @[:@524.4]
  output         io_inst_st_valid, // @[:@524.4]
  output [127:0] io_inst_st_bits // @[:@524.4]
);
  wire  inst_q_clock; // @[Fetch.scala 57:22:@526.4]
  wire  inst_q_reset; // @[Fetch.scala 57:22:@526.4]
  wire  inst_q_io_enq_ready; // @[Fetch.scala 57:22:@526.4]
  wire  inst_q_io_enq_valid; // @[Fetch.scala 57:22:@526.4]
  wire [127:0] inst_q_io_enq_bits; // @[Fetch.scala 57:22:@526.4]
  wire  inst_q_io_deq_ready; // @[Fetch.scala 57:22:@526.4]
  wire  inst_q_io_deq_valid; // @[Fetch.scala 57:22:@526.4]
  wire [127:0] inst_q_io_deq_bits; // @[Fetch.scala 57:22:@526.4]
  wire [7:0] inst_q_io_count; // @[Fetch.scala 57:22:@526.4]
  wire [127:0] dec_io_inst; // @[Fetch.scala 58:19:@529.4]
  wire  dec_io_isLoad; // @[Fetch.scala 58:19:@529.4]
  wire  dec_io_isCompute; // @[Fetch.scala 58:19:@529.4]
  wire  dec_io_isStore; // @[Fetch.scala 58:19:@529.4]
  reg  s1_launch; // @[Fetch.scala 60:26:@532.4]
  reg [31:0] _RAND_0;
  wire  _T_65; // @[Fetch.scala 61:27:@534.4]
  wire  pulse; // @[Fetch.scala 61:25:@535.4]
  reg [31:0] raddr; // @[Fetch.scala 63:18:@536.4]
  reg [31:0] _RAND_1;
  reg [7:0] rlen; // @[Fetch.scala 64:17:@537.4]
  reg [31:0] _RAND_2;
  reg [7:0] ilen; // @[Fetch.scala 65:17:@538.4]
  reg [31:0] _RAND_3;
  reg [31:0] xrem; // @[Fetch.scala 67:17:@539.4]
  reg [31:0] _RAND_4;
  wire [32:0] _GEN_46; // @[Fetch.scala 68:29:@540.4]
  wire [32:0] _T_71; // @[Fetch.scala 68:29:@540.4]
  wire [33:0] _T_73; // @[Fetch.scala 68:37:@541.4]
  wire [33:0] _T_74; // @[Fetch.scala 68:37:@542.4]
  wire [32:0] xsize; // @[Fetch.scala 68:37:@543.4]
  reg [2:0] state; // @[Fetch.scala 73:22:@544.4]
  reg [31:0] _RAND_5;
  wire  _T_76; // @[Conditional.scala 37:30:@545.4]
  wire  _T_77; // @[Fetch.scala 80:20:@549.8]
  wire [32:0] _T_79; // @[Fetch.scala 82:25:@552.10]
  wire [9:0] _T_82; // @[Fetch.scala 85:24:@557.10]
  wire [9:0] _T_83; // @[Fetch.scala 85:24:@558.10]
  wire [8:0] _T_84; // @[Fetch.scala 85:24:@559.10]
  wire [8:0] _T_86; // @[Fetch.scala 86:25:@561.10]
  wire [9:0] _T_88; // @[Fetch.scala 86:33:@562.10]
  wire [9:0] _T_89; // @[Fetch.scala 86:33:@563.10]
  wire [8:0] _T_90; // @[Fetch.scala 86:33:@564.10]
  wire [33:0] _T_91; // @[Fetch.scala 87:25:@566.10]
  wire [33:0] _T_92; // @[Fetch.scala 87:25:@567.10]
  wire [32:0] _T_93; // @[Fetch.scala 87:25:@568.10]
  wire [32:0] _GEN_0; // @[Fetch.scala 80:28:@550.8]
  wire [32:0] _GEN_1; // @[Fetch.scala 80:28:@550.8]
  wire [32:0] _GEN_2; // @[Fetch.scala 80:28:@550.8]
  wire [2:0] _GEN_3; // @[Fetch.scala 78:19:@547.6]
  wire [32:0] _GEN_4; // @[Fetch.scala 78:19:@547.6]
  wire [32:0] _GEN_5; // @[Fetch.scala 78:19:@547.6]
  wire [32:0] _GEN_6; // @[Fetch.scala 78:19:@547.6]
  wire  _T_94; // @[Conditional.scala 37:30:@574.6]
  wire [2:0] _GEN_7; // @[Fetch.scala 92:33:@576.8]
  wire  _T_95; // @[Conditional.scala 37:30:@581.8]
  wire [2:0] _GEN_8; // @[Fetch.scala 97:34:@583.10]
  wire  _T_96; // @[Conditional.scala 37:30:@588.10]
  wire  _T_97; // @[Fetch.scala 103:30:@591.14]
  wire [2:0] _GEN_9; // @[Fetch.scala 103:40:@592.14]
  wire [2:0] _GEN_10; // @[Fetch.scala 102:34:@590.12]
  wire  _T_98; // @[Conditional.scala 37:30:@601.12]
  wire  _T_100; // @[Fetch.scala 111:28:@603.14]
  wire  _T_102; // @[Fetch.scala 112:19:@605.16]
  wire  _T_103; // @[Fetch.scala 114:25:@610.18]
  wire [31:0] _T_105; // @[Fetch.scala 117:24:@614.20]
  wire [32:0] _T_117; // @[Fetch.scala 123:24:@629.20]
  wire [32:0] _T_118; // @[Fetch.scala 123:24:@630.20]
  wire [31:0] _T_119; // @[Fetch.scala 123:24:@631.20]
  wire [31:0] _GEN_12; // @[Fetch.scala 114:33:@611.18]
  wire [31:0] _GEN_13; // @[Fetch.scala 114:33:@611.18]
  wire [31:0] _GEN_14; // @[Fetch.scala 114:33:@611.18]
  wire [2:0] _GEN_15; // @[Fetch.scala 112:28:@606.16]
  wire [31:0] _GEN_16; // @[Fetch.scala 112:28:@606.16]
  wire [31:0] _GEN_17; // @[Fetch.scala 112:28:@606.16]
  wire [31:0] _GEN_18; // @[Fetch.scala 112:28:@606.16]
  wire [2:0] _GEN_19; // @[Fetch.scala 111:37:@604.14]
  wire [31:0] _GEN_20; // @[Fetch.scala 111:37:@604.14]
  wire [31:0] _GEN_21; // @[Fetch.scala 111:37:@604.14]
  wire [31:0] _GEN_22; // @[Fetch.scala 111:37:@604.14]
  wire [2:0] _GEN_23; // @[Conditional.scala 39:67:@602.12]
  wire [31:0] _GEN_24; // @[Conditional.scala 39:67:@602.12]
  wire [31:0] _GEN_25; // @[Conditional.scala 39:67:@602.12]
  wire [31:0] _GEN_26; // @[Conditional.scala 39:67:@602.12]
  wire [2:0] _GEN_27; // @[Conditional.scala 39:67:@589.10]
  wire [31:0] _GEN_28; // @[Conditional.scala 39:67:@589.10]
  wire [31:0] _GEN_29; // @[Conditional.scala 39:67:@589.10]
  wire [31:0] _GEN_30; // @[Conditional.scala 39:67:@589.10]
  wire [2:0] _GEN_31; // @[Conditional.scala 39:67:@582.8]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67:@582.8]
  wire [31:0] _GEN_33; // @[Conditional.scala 39:67:@582.8]
  wire [31:0] _GEN_34; // @[Conditional.scala 39:67:@582.8]
  wire [2:0] _GEN_35; // @[Conditional.scala 39:67:@575.6]
  wire [31:0] _GEN_36; // @[Conditional.scala 39:67:@575.6]
  wire [31:0] _GEN_37; // @[Conditional.scala 39:67:@575.6]
  wire [31:0] _GEN_38; // @[Conditional.scala 39:67:@575.6]
  wire [2:0] _GEN_39; // @[Conditional.scala 40:58:@546.4]
  wire [32:0] _GEN_40; // @[Conditional.scala 40:58:@546.4]
  wire [32:0] _GEN_41; // @[Conditional.scala 40:58:@546.4]
  wire [32:0] _GEN_42; // @[Conditional.scala 40:58:@546.4]
  wire  _T_120; // @[Fetch.scala 130:14:@636.4]
  wire  _T_121; // @[Fetch.scala 132:20:@641.6]
  wire  _T_124; // @[Fetch.scala 132:31:@643.6]
  wire  _T_126; // @[Fetch.scala 132:66:@644.6]
  wire  _T_127; // @[Fetch.scala 132:58:@645.6]
  wire [32:0] _T_128; // @[Fetch.scala 133:20:@647.8]
  wire [31:0] _T_129; // @[Fetch.scala 133:20:@648.8]
  wire [31:0] _GEN_43; // @[Fetch.scala 132:75:@646.6]
  reg [63:0] lsb; // @[Fetch.scala 142:16:@656.4]
  reg [63:0] _RAND_6;
  wire  _T_132; // @[Fetch.scala 146:14:@658.4]
  wire  _T_133; // @[Fetch.scala 148:55:@662.4]
  wire  _T_135; // @[Fetch.scala 155:37:@667.4]
  wire  _T_138; // @[Fetch.scala 156:40:@671.4]
  wire  _T_141; // @[Fetch.scala 157:38:@675.4]
  wire [2:0] deq_sel; // @[Cat.scala 30:58:@683.4]
  wire  _T_149; // @[Mux.scala 46:19:@684.4]
  wire  _T_150; // @[Mux.scala 46:16:@685.4]
  wire  _T_151; // @[Mux.scala 46:19:@686.4]
  wire  _T_152; // @[Mux.scala 46:16:@687.4]
  wire  _T_153; // @[Mux.scala 46:19:@688.4]
  wire  deq_ready; // @[Mux.scala 46:16:@689.4]
  wire  _T_154; // @[Fetch.scala 175:36:@690.4]
  Queue inst_q ( // @[Fetch.scala 57:22:@526.4]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits),
    .io_count(inst_q_io_count)
  );
  FetchDecode dec ( // @[Fetch.scala 58:19:@529.4]
    .io_inst(dec_io_inst),
    .io_isLoad(dec_io_isLoad),
    .io_isCompute(dec_io_isCompute),
    .io_isStore(dec_io_isStore)
  );
  assign _T_65 = ~ s1_launch; // @[Fetch.scala 61:27:@534.4]
  assign pulse = io_launch & _T_65; // @[Fetch.scala 61:25:@535.4]
  assign _GEN_46 = {{1'd0}, io_ins_count}; // @[Fetch.scala 68:29:@540.4]
  assign _T_71 = _GEN_46 << 1'h1; // @[Fetch.scala 68:29:@540.4]
  assign _T_73 = _T_71 - 33'h1; // @[Fetch.scala 68:37:@541.4]
  assign _T_74 = $unsigned(_T_73); // @[Fetch.scala 68:37:@542.4]
  assign xsize = _T_74[32:0]; // @[Fetch.scala 68:37:@543.4]
  assign _T_76 = 3'h0 == state; // @[Conditional.scala 37:30:@545.4]
  assign _T_77 = xsize < 33'h100; // @[Fetch.scala 80:20:@549.8]
  assign _T_79 = xsize >> 1'h1; // @[Fetch.scala 82:25:@552.10]
  assign _T_82 = 9'h100 - 9'h1; // @[Fetch.scala 85:24:@557.10]
  assign _T_83 = $unsigned(_T_82); // @[Fetch.scala 85:24:@558.10]
  assign _T_84 = _T_83[8:0]; // @[Fetch.scala 85:24:@559.10]
  assign _T_86 = 9'h100 >> 1'h1; // @[Fetch.scala 86:25:@561.10]
  assign _T_88 = _T_86 - 9'h1; // @[Fetch.scala 86:33:@562.10]
  assign _T_89 = $unsigned(_T_88); // @[Fetch.scala 86:33:@563.10]
  assign _T_90 = _T_89[8:0]; // @[Fetch.scala 86:33:@564.10]
  assign _T_91 = xsize - 33'h100; // @[Fetch.scala 87:25:@566.10]
  assign _T_92 = $unsigned(_T_91); // @[Fetch.scala 87:25:@567.10]
  assign _T_93 = _T_92[32:0]; // @[Fetch.scala 87:25:@568.10]
  assign _GEN_0 = _T_77 ? xsize : {{24'd0}, _T_84}; // @[Fetch.scala 80:28:@550.8]
  assign _GEN_1 = _T_77 ? _T_79 : {{24'd0}, _T_90}; // @[Fetch.scala 80:28:@550.8]
  assign _GEN_2 = _T_77 ? 33'h0 : _T_93; // @[Fetch.scala 80:28:@550.8]
  assign _GEN_3 = pulse ? 3'h1 : state; // @[Fetch.scala 78:19:@547.6]
  assign _GEN_4 = pulse ? _GEN_0 : {{25'd0}, rlen}; // @[Fetch.scala 78:19:@547.6]
  assign _GEN_5 = pulse ? _GEN_1 : {{25'd0}, ilen}; // @[Fetch.scala 78:19:@547.6]
  assign _GEN_6 = pulse ? _GEN_2 : {{1'd0}, xrem}; // @[Fetch.scala 78:19:@547.6]
  assign _T_94 = 3'h1 == state; // @[Conditional.scala 37:30:@574.6]
  assign _GEN_7 = io_vme_rd_cmd_ready ? 3'h2 : state; // @[Fetch.scala 92:33:@576.8]
  assign _T_95 = 3'h2 == state; // @[Conditional.scala 37:30:@581.8]
  assign _GEN_8 = io_vme_rd_data_valid ? 3'h3 : state; // @[Fetch.scala 97:34:@583.10]
  assign _T_96 = 3'h3 == state; // @[Conditional.scala 37:30:@588.10]
  assign _T_97 = inst_q_io_count == ilen; // @[Fetch.scala 103:30:@591.14]
  assign _GEN_9 = _T_97 ? 3'h4 : 3'h2; // @[Fetch.scala 103:40:@592.14]
  assign _GEN_10 = io_vme_rd_data_valid ? _GEN_9 : state; // @[Fetch.scala 102:34:@590.12]
  assign _T_98 = 3'h4 == state; // @[Conditional.scala 37:30:@601.12]
  assign _T_100 = inst_q_io_count == 8'h0; // @[Fetch.scala 111:28:@603.14]
  assign _T_102 = xrem == 32'h0; // @[Fetch.scala 112:19:@605.16]
  assign _T_103 = xrem < 32'h100; // @[Fetch.scala 114:25:@610.18]
  assign _T_105 = xrem >> 1'h1; // @[Fetch.scala 117:24:@614.20]
  assign _T_117 = xrem - 32'h100; // @[Fetch.scala 123:24:@629.20]
  assign _T_118 = $unsigned(_T_117); // @[Fetch.scala 123:24:@630.20]
  assign _T_119 = _T_118[31:0]; // @[Fetch.scala 123:24:@631.20]
  assign _GEN_12 = _T_103 ? xrem : {{23'd0}, _T_84}; // @[Fetch.scala 114:33:@611.18]
  assign _GEN_13 = _T_103 ? _T_105 : {{23'd0}, _T_90}; // @[Fetch.scala 114:33:@611.18]
  assign _GEN_14 = _T_103 ? 32'h0 : _T_119; // @[Fetch.scala 114:33:@611.18]
  assign _GEN_15 = _T_102 ? 3'h0 : 3'h1; // @[Fetch.scala 112:28:@606.16]
  assign _GEN_16 = _T_102 ? {{24'd0}, rlen} : _GEN_12; // @[Fetch.scala 112:28:@606.16]
  assign _GEN_17 = _T_102 ? {{24'd0}, ilen} : _GEN_13; // @[Fetch.scala 112:28:@606.16]
  assign _GEN_18 = _T_102 ? xrem : _GEN_14; // @[Fetch.scala 112:28:@606.16]
  assign _GEN_19 = _T_100 ? _GEN_15 : state; // @[Fetch.scala 111:37:@604.14]
  assign _GEN_20 = _T_100 ? _GEN_16 : {{24'd0}, rlen}; // @[Fetch.scala 111:37:@604.14]
  assign _GEN_21 = _T_100 ? _GEN_17 : {{24'd0}, ilen}; // @[Fetch.scala 111:37:@604.14]
  assign _GEN_22 = _T_100 ? _GEN_18 : xrem; // @[Fetch.scala 111:37:@604.14]
  assign _GEN_23 = _T_98 ? _GEN_19 : state; // @[Conditional.scala 39:67:@602.12]
  assign _GEN_24 = _T_98 ? _GEN_20 : {{24'd0}, rlen}; // @[Conditional.scala 39:67:@602.12]
  assign _GEN_25 = _T_98 ? _GEN_21 : {{24'd0}, ilen}; // @[Conditional.scala 39:67:@602.12]
  assign _GEN_26 = _T_98 ? _GEN_22 : xrem; // @[Conditional.scala 39:67:@602.12]
  assign _GEN_27 = _T_96 ? _GEN_10 : _GEN_23; // @[Conditional.scala 39:67:@589.10]
  assign _GEN_28 = _T_96 ? {{24'd0}, rlen} : _GEN_24; // @[Conditional.scala 39:67:@589.10]
  assign _GEN_29 = _T_96 ? {{24'd0}, ilen} : _GEN_25; // @[Conditional.scala 39:67:@589.10]
  assign _GEN_30 = _T_96 ? xrem : _GEN_26; // @[Conditional.scala 39:67:@589.10]
  assign _GEN_31 = _T_95 ? _GEN_8 : _GEN_27; // @[Conditional.scala 39:67:@582.8]
  assign _GEN_32 = _T_95 ? {{24'd0}, rlen} : _GEN_28; // @[Conditional.scala 39:67:@582.8]
  assign _GEN_33 = _T_95 ? {{24'd0}, ilen} : _GEN_29; // @[Conditional.scala 39:67:@582.8]
  assign _GEN_34 = _T_95 ? xrem : _GEN_30; // @[Conditional.scala 39:67:@582.8]
  assign _GEN_35 = _T_94 ? _GEN_7 : _GEN_31; // @[Conditional.scala 39:67:@575.6]
  assign _GEN_36 = _T_94 ? {{24'd0}, rlen} : _GEN_32; // @[Conditional.scala 39:67:@575.6]
  assign _GEN_37 = _T_94 ? {{24'd0}, ilen} : _GEN_33; // @[Conditional.scala 39:67:@575.6]
  assign _GEN_38 = _T_94 ? xrem : _GEN_34; // @[Conditional.scala 39:67:@575.6]
  assign _GEN_39 = _T_76 ? _GEN_3 : _GEN_35; // @[Conditional.scala 40:58:@546.4]
  assign _GEN_40 = _T_76 ? _GEN_4 : {{1'd0}, _GEN_36}; // @[Conditional.scala 40:58:@546.4]
  assign _GEN_41 = _T_76 ? _GEN_5 : {{1'd0}, _GEN_37}; // @[Conditional.scala 40:58:@546.4]
  assign _GEN_42 = _T_76 ? _GEN_6 : {{1'd0}, _GEN_38}; // @[Conditional.scala 40:58:@546.4]
  assign _T_120 = state == 3'h0; // @[Fetch.scala 130:14:@636.4]
  assign _T_121 = state == 3'h4; // @[Fetch.scala 132:20:@641.6]
  assign _T_124 = _T_121 & _T_100; // @[Fetch.scala 132:31:@643.6]
  assign _T_126 = xrem != 32'h0; // @[Fetch.scala 132:66:@644.6]
  assign _T_127 = _T_124 & _T_126; // @[Fetch.scala 132:58:@645.6]
  assign _T_128 = raddr + 32'h800; // @[Fetch.scala 133:20:@647.8]
  assign _T_129 = raddr + 32'h800; // @[Fetch.scala 133:20:@648.8]
  assign _GEN_43 = _T_127 ? _T_129 : raddr; // @[Fetch.scala 132:75:@646.6]
  assign _T_132 = state == 3'h2; // @[Fetch.scala 146:14:@658.4]
  assign _T_133 = state == 3'h3; // @[Fetch.scala 148:55:@662.4]
  assign _T_135 = dec_io_isLoad & inst_q_io_deq_valid; // @[Fetch.scala 155:37:@667.4]
  assign _T_138 = dec_io_isCompute & inst_q_io_deq_valid; // @[Fetch.scala 156:40:@671.4]
  assign _T_141 = dec_io_isStore & inst_q_io_deq_valid; // @[Fetch.scala 157:38:@675.4]
  assign deq_sel = {dec_io_isCompute,dec_io_isStore,dec_io_isLoad}; // @[Cat.scala 30:58:@683.4]
  assign _T_149 = 3'h4 == deq_sel; // @[Mux.scala 46:19:@684.4]
  assign _T_150 = _T_149 ? io_inst_co_ready : 1'h0; // @[Mux.scala 46:16:@685.4]
  assign _T_151 = 3'h2 == deq_sel; // @[Mux.scala 46:19:@686.4]
  assign _T_152 = _T_151 ? io_inst_st_ready : _T_150; // @[Mux.scala 46:16:@687.4]
  assign _T_153 = 3'h1 == deq_sel; // @[Mux.scala 46:19:@688.4]
  assign deq_ready = _T_153 ? io_inst_ld_ready : _T_152; // @[Mux.scala 46:16:@689.4]
  assign _T_154 = deq_ready & inst_q_io_deq_valid; // @[Fetch.scala 175:36:@690.4]
  assign io_vme_rd_cmd_valid = state == 3'h1; // @[Fetch.scala 136:23:@652.4]
  assign io_vme_rd_cmd_bits_addr = raddr; // @[Fetch.scala 137:27:@653.4]
  assign io_vme_rd_cmd_bits_len = rlen; // @[Fetch.scala 138:26:@654.4]
  assign io_vme_rd_data_ready = inst_q_io_enq_ready; // @[Fetch.scala 140:24:@655.4]
  assign io_inst_ld_valid = _T_135 & _T_121; // @[Fetch.scala 155:20:@670.4]
  assign io_inst_ld_bits = inst_q_io_deq_bits; // @[Fetch.scala 159:19:@679.4]
  assign io_inst_co_valid = _T_138 & _T_121; // @[Fetch.scala 156:20:@674.4]
  assign io_inst_co_bits = inst_q_io_deq_bits; // @[Fetch.scala 160:19:@680.4]
  assign io_inst_st_valid = _T_141 & _T_121; // @[Fetch.scala 157:20:@678.4]
  assign io_inst_st_bits = inst_q_io_deq_bits; // @[Fetch.scala 161:19:@681.4]
  assign inst_q_clock = clock; // @[:@527.4]
  assign inst_q_reset = reset; // @[:@528.4]
  assign inst_q_io_enq_valid = io_vme_rd_data_valid & _T_133; // @[Fetch.scala 148:23:@664.4]
  assign inst_q_io_enq_bits = {io_vme_rd_data_bits,lsb}; // @[Fetch.scala 149:22:@665.4]
  assign inst_q_io_deq_ready = _T_154 & _T_121; // @[Fetch.scala 175:23:@693.4]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Fetch.scala 152:15:@666.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_launch = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  raddr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rlen = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ilen = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xrem = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{`RANDOM}};
  lsb = _RAND_6[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    s1_launch <= io_launch;
    if (_T_120) begin
      raddr <= io_ins_baddr;
    end else begin
      if (_T_127) begin
        raddr <= _T_129;
      end
    end
    rlen <= _GEN_40[7:0];
    ilen <= _GEN_41[7:0];
    xrem <= _GEN_42[31:0];
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_76) begin
        if (pulse) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_94) begin
          if (io_vme_rd_cmd_ready) begin
            state <= 3'h2;
          end
        end else begin
          if (_T_95) begin
            if (io_vme_rd_data_valid) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_96) begin
              if (io_vme_rd_data_valid) begin
                if (_T_97) begin
                  state <= 3'h4;
                end else begin
                  state <= 3'h2;
                end
              end
            end else begin
              if (_T_98) begin
                if (_T_100) begin
                  if (_T_102) begin
                    state <= 3'h0;
                  end else begin
                    state <= 3'h1;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_132) begin
      lsb <= io_vme_rd_data_bits;
    end
  end
endmodule
module Semaphore( // @[:@695.2]
  input   clock, // @[:@696.4]
  input   reset, // @[:@697.4]
  input   io_spost, // @[:@698.4]
  input   io_swait, // @[:@698.4]
  output  io_sready // @[:@698.4]
);
  reg [7:0] cnt; // @[Semaphore.scala 38:20:@700.4]
  reg [31:0] _RAND_0;
  wire  _T_14; // @[Semaphore.scala 39:20:@701.4]
  wire  _T_15; // @[Semaphore.scala 39:17:@702.4]
  wire  _T_17; // @[Semaphore.scala 39:37:@703.4]
  wire  _T_18; // @[Semaphore.scala 39:30:@704.4]
  wire [8:0] _T_20; // @[Semaphore.scala 40:16:@706.6]
  wire [7:0] _T_21; // @[Semaphore.scala 40:16:@707.6]
  wire [7:0] _GEN_0; // @[Semaphore.scala 39:74:@705.4]
  wire  _T_23; // @[Semaphore.scala 42:8:@710.4]
  wire  _T_24; // @[Semaphore.scala 42:18:@711.4]
  wire  _T_26; // @[Semaphore.scala 42:37:@712.4]
  wire  _T_27; // @[Semaphore.scala 42:30:@713.4]
  wire [8:0] _T_29; // @[Semaphore.scala 42:59:@715.6]
  wire [8:0] _T_30; // @[Semaphore.scala 42:59:@716.6]
  wire [7:0] _T_31; // @[Semaphore.scala 42:59:@717.6]
  wire [7:0] _GEN_1; // @[Semaphore.scala 42:46:@714.4]
  assign _T_14 = io_swait == 1'h0; // @[Semaphore.scala 39:20:@701.4]
  assign _T_15 = io_spost & _T_14; // @[Semaphore.scala 39:17:@702.4]
  assign _T_17 = cnt != 8'hff; // @[Semaphore.scala 39:37:@703.4]
  assign _T_18 = _T_15 & _T_17; // @[Semaphore.scala 39:30:@704.4]
  assign _T_20 = cnt + 8'h1; // @[Semaphore.scala 40:16:@706.6]
  assign _T_21 = cnt + 8'h1; // @[Semaphore.scala 40:16:@707.6]
  assign _GEN_0 = _T_18 ? _T_21 : cnt; // @[Semaphore.scala 39:74:@705.4]
  assign _T_23 = io_spost == 1'h0; // @[Semaphore.scala 42:8:@710.4]
  assign _T_24 = _T_23 & io_swait; // @[Semaphore.scala 42:18:@711.4]
  assign _T_26 = cnt != 8'h0; // @[Semaphore.scala 42:37:@712.4]
  assign _T_27 = _T_24 & _T_26; // @[Semaphore.scala 42:30:@713.4]
  assign _T_29 = cnt - 8'h1; // @[Semaphore.scala 42:59:@715.6]
  assign _T_30 = $unsigned(_T_29); // @[Semaphore.scala 42:59:@716.6]
  assign _T_31 = _T_30[7:0]; // @[Semaphore.scala 42:59:@717.6]
  assign _GEN_1 = _T_27 ? _T_31 : _GEN_0; // @[Semaphore.scala 42:46:@714.4]
  assign io_sready = cnt != 8'h0; // @[Semaphore.scala 43:13:@721.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 8'h0;
    end else begin
      if (_T_27) begin
        cnt <= _T_31;
      end else begin
        if (_T_18) begin
          cnt <= _T_21;
        end
      end
    end
  end
endmodule
module Queue_1( // @[:@723.2]
  input          clock, // @[:@724.4]
  input          reset, // @[:@725.4]
  output         io_enq_ready, // @[:@726.4]
  input          io_enq_valid, // @[:@726.4]
  input  [127:0] io_enq_bits, // @[:@726.4]
  input          io_deq_ready, // @[:@726.4]
  output         io_deq_valid, // @[:@726.4]
  output [127:0] io_deq_bits // @[:@726.4]
);
  reg [127:0] _T_35 [0:511]; // @[Decoupled.scala 215:24:@728.4]
  reg [127:0] _RAND_0;
  wire [127:0] _T_35__T_68_data; // @[Decoupled.scala 215:24:@728.4]
  wire [8:0] _T_35__T_68_addr; // @[Decoupled.scala 215:24:@728.4]
  wire [127:0] _T_35__T_54_data; // @[Decoupled.scala 215:24:@728.4]
  wire [8:0] _T_35__T_54_addr; // @[Decoupled.scala 215:24:@728.4]
  wire  _T_35__T_54_mask; // @[Decoupled.scala 215:24:@728.4]
  wire  _T_35__T_54_en; // @[Decoupled.scala 215:24:@728.4]
  reg [8:0] value; // @[Counter.scala 26:33:@729.4]
  reg [31:0] _RAND_1;
  reg [8:0] value_1; // @[Counter.scala 26:33:@730.4]
  reg [31:0] _RAND_2;
  reg  _T_42; // @[Decoupled.scala 218:35:@731.4]
  reg [31:0] _RAND_3;
  wire  _T_43; // @[Decoupled.scala 220:41:@732.4]
  wire  _T_45; // @[Decoupled.scala 221:36:@733.4]
  wire  _T_46; // @[Decoupled.scala 221:33:@734.4]
  wire  _T_47; // @[Decoupled.scala 222:32:@735.4]
  wire  _T_48; // @[Decoupled.scala 37:37:@736.4]
  wire  _T_51; // @[Decoupled.scala 37:37:@739.4]
  wire [9:0] _T_57; // @[Counter.scala 35:22:@746.6]
  wire [8:0] _T_58; // @[Counter.scala 35:22:@747.6]
  wire [8:0] _GEN_5; // @[Decoupled.scala 226:17:@742.4]
  wire [9:0] _T_61; // @[Counter.scala 35:22:@752.6]
  wire [8:0] _T_62; // @[Counter.scala 35:22:@753.6]
  wire [8:0] _GEN_6; // @[Decoupled.scala 230:17:@750.4]
  wire  _T_63; // @[Decoupled.scala 233:16:@756.4]
  wire  _GEN_7; // @[Decoupled.scala 233:28:@757.4]
  assign _T_35__T_68_addr = value_1;
  assign _T_35__T_68_data = _T_35[_T_35__T_68_addr]; // @[Decoupled.scala 215:24:@728.4]
  assign _T_35__T_54_data = io_enq_bits;
  assign _T_35__T_54_addr = value;
  assign _T_35__T_54_mask = 1'h1;
  assign _T_35__T_54_en = io_enq_ready & io_enq_valid;
  assign _T_43 = value == value_1; // @[Decoupled.scala 220:41:@732.4]
  assign _T_45 = _T_42 == 1'h0; // @[Decoupled.scala 221:36:@733.4]
  assign _T_46 = _T_43 & _T_45; // @[Decoupled.scala 221:33:@734.4]
  assign _T_47 = _T_43 & _T_42; // @[Decoupled.scala 222:32:@735.4]
  assign _T_48 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:@736.4]
  assign _T_51 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:@739.4]
  assign _T_57 = value + 9'h1; // @[Counter.scala 35:22:@746.6]
  assign _T_58 = value + 9'h1; // @[Counter.scala 35:22:@747.6]
  assign _GEN_5 = _T_48 ? _T_58 : value; // @[Decoupled.scala 226:17:@742.4]
  assign _T_61 = value_1 + 9'h1; // @[Counter.scala 35:22:@752.6]
  assign _T_62 = value_1 + 9'h1; // @[Counter.scala 35:22:@753.6]
  assign _GEN_6 = _T_51 ? _T_62 : value_1; // @[Decoupled.scala 230:17:@750.4]
  assign _T_63 = _T_48 != _T_51; // @[Decoupled.scala 233:16:@756.4]
  assign _GEN_7 = _T_63 ? _T_48 : _T_42; // @[Decoupled.scala 233:28:@757.4]
  assign io_enq_ready = _T_47 == 1'h0; // @[Decoupled.scala 238:16:@763.4]
  assign io_deq_valid = _T_46 == 1'h0; // @[Decoupled.scala 237:16:@761.4]
  assign io_deq_bits = _T_35__T_68_data; // @[Decoupled.scala 239:15:@765.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    _T_35[initvar] = _RAND_0[127:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_42 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35__T_54_en & _T_35__T_54_mask) begin
      _T_35[_T_35__T_54_addr] <= _T_35__T_54_data; // @[Decoupled.scala 215:24:@728.4]
    end
    if (reset) begin
      value <= 9'h0;
    end else begin
      if (_T_48) begin
        value <= _T_58;
      end
    end
    if (reset) begin
      value_1 <= 9'h0;
    end else begin
      if (_T_51) begin
        value_1 <= _T_62;
      end
    end
    if (reset) begin
      _T_42 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_42 <= _T_48;
      end
    end
  end
endmodule
module LoadDecode( // @[:@774.2]
  input  [127:0] io_inst, // @[:@777.4]
  output         io_push_next, // @[:@777.4]
  output         io_pop_next, // @[:@777.4]
  output         io_isInput, // @[:@777.4]
  output         io_isWeight, // @[:@777.4]
  output         io_isSync // @[:@777.4]
);
  wire [15:0] dec_xsize; // @[Decode.scala 174:29:@802.4]
  wire [127:0] _T_39; // @[Decode.scala 177:25:@816.4]
  wire  _T_40; // @[Decode.scala 177:25:@817.4]
  wire  _T_42; // @[Decode.scala 177:46:@818.4]
  wire  _T_47; // @[Decode.scala 178:26:@822.4]
  wire  _T_59; // @[Decode.scala 179:34:@830.4]
  wire  _T_61; // @[Decode.scala 179:66:@831.4]
  assign dec_xsize = io_inst[95:80]; // @[Decode.scala 174:29:@802.4]
  assign _T_39 = io_inst & 128'h187; // @[Decode.scala 177:25:@816.4]
  assign _T_40 = 128'h100 == _T_39; // @[Decode.scala 177:25:@817.4]
  assign _T_42 = dec_xsize != 16'h0; // @[Decode.scala 177:46:@818.4]
  assign _T_47 = 128'h80 == _T_39; // @[Decode.scala 178:26:@822.4]
  assign _T_59 = _T_40 | _T_47; // @[Decode.scala 179:34:@830.4]
  assign _T_61 = dec_xsize == 16'h0; // @[Decode.scala 179:66:@831.4]
  assign io_push_next = io_inst[6]; // @[Decode.scala 175:16:@814.4]
  assign io_pop_next = io_inst[4]; // @[Decode.scala 176:15:@815.4]
  assign io_isInput = _T_40 & _T_42; // @[Decode.scala 177:14:@820.4]
  assign io_isWeight = _T_47 & _T_42; // @[Decode.scala 178:15:@825.4]
  assign io_isSync = _T_59 & _T_61; // @[Decode.scala 179:13:@833.4]
endmodule
module TensorDataCtrl( // @[:@835.2]
  input          clock, // @[:@836.4]
  input          io_start, // @[:@838.4]
  output         io_done, // @[:@838.4]
  input  [127:0] io_inst, // @[:@838.4]
  input  [31:0]  io_baddr, // @[:@838.4]
  input          io_xinit, // @[:@838.4]
  input          io_xupdate, // @[:@838.4]
  input          io_yupdate, // @[:@838.4]
  output         io_stride, // @[:@838.4]
  output         io_split, // @[:@838.4]
  output [31:0]  io_addr, // @[:@838.4]
  output [7:0]   io_len // @[:@838.4]
);
  wire [31:0] dec_dram_offset; // @[TensorUtil.scala 251:29:@857.4]
  wire [15:0] dec_ysize; // @[TensorUtil.scala 251:29:@861.4]
  wire [15:0] dec_xsize; // @[TensorUtil.scala 251:29:@863.4]
  wire [15:0] dec_xstride; // @[TensorUtil.scala 251:29:@865.4]
  reg [31:0] caddr; // @[TensorUtil.scala 253:18:@875.4]
  reg [31:0] _RAND_0;
  reg [31:0] baddr; // @[TensorUtil.scala 254:18:@876.4]
  reg [31:0] _RAND_1;
  reg [7:0] len; // @[TensorUtil.scala 255:16:@877.4]
  reg [31:0] _RAND_2;
  reg [7:0] xcnt; // @[TensorUtil.scala 267:17:@942.4]
  reg [31:0] _RAND_3;
  reg [15:0] xrem; // @[TensorUtil.scala 268:17:@943.4]
  reg [31:0] _RAND_4;
  wire [16:0] _GEN_27; // @[TensorUtil.scala 269:26:@944.4]
  wire [16:0] _T_154; // @[TensorUtil.scala 269:26:@944.4]
  wire [17:0] _T_156; // @[TensorUtil.scala 269:51:@945.4]
  wire [17:0] _T_157; // @[TensorUtil.scala 269:51:@946.4]
  wire [16:0] xsize; // @[TensorUtil.scala 269:51:@947.4]
  reg [15:0] ycnt; // @[TensorUtil.scala 271:17:@948.4]
  reg [31:0] _RAND_5;
  reg [31:0] xfer_bytes; // @[TensorUtil.scala 273:23:@949.4]
  reg [31:0] _RAND_6;
  wire [19:0] _GEN_28; // @[TensorUtil.scala 275:35:@950.4]
  wire [19:0] xstride_bytes; // @[TensorUtil.scala 275:35:@950.4]
  wire [35:0] _GEN_29; // @[TensorUtil.scala 277:66:@951.4]
  wire [35:0] _T_160; // @[TensorUtil.scala 277:66:@951.4]
  wire [35:0] _T_161; // @[TensorUtil.scala 277:47:@952.4]
  wire [35:0] _GEN_30; // @[TensorUtil.scala 277:33:@953.4]
  wire [35:0] xfer_init_addr; // @[TensorUtil.scala 277:33:@953.4]
  wire [32:0] _T_162; // @[TensorUtil.scala 278:31:@954.4]
  wire [31:0] xfer_split_addr; // @[TensorUtil.scala 278:31:@955.4]
  wire [31:0] _GEN_31; // @[TensorUtil.scala 279:32:@956.4]
  wire [32:0] _T_163; // @[TensorUtil.scala 279:32:@956.4]
  wire [31:0] xfer_stride_addr; // @[TensorUtil.scala 279:32:@957.4]
  wire [35:0] _GEN_12; // @[TensorUtil.scala 281:55:@958.4]
  wire [11:0] _T_164; // @[TensorUtil.scala 281:55:@958.4]
  wire [12:0] _T_165; // @[TensorUtil.scala 281:38:@959.4]
  wire [12:0] _T_166; // @[TensorUtil.scala 281:38:@960.4]
  wire [11:0] xfer_init_bytes; // @[TensorUtil.scala 281:38:@961.4]
  wire [8:0] xfer_init_pulses; // @[TensorUtil.scala 282:43:@962.4]
  wire [31:0] _GEN_16; // @[TensorUtil.scala 283:56:@963.4]
  wire [11:0] _T_167; // @[TensorUtil.scala 283:56:@963.4]
  wire [12:0] _T_168; // @[TensorUtil.scala 283:38:@964.4]
  wire [12:0] _T_169; // @[TensorUtil.scala 283:38:@965.4]
  wire [11:0] xfer_split_bytes; // @[TensorUtil.scala 283:38:@966.4]
  wire [8:0] xfer_split_pulses; // @[TensorUtil.scala 284:44:@967.4]
  wire [31:0] _GEN_18; // @[TensorUtil.scala 285:57:@968.4]
  wire [11:0] _T_170; // @[TensorUtil.scala 285:57:@968.4]
  wire [12:0] _T_171; // @[TensorUtil.scala 285:38:@969.4]
  wire [12:0] _T_172; // @[TensorUtil.scala 285:38:@970.4]
  wire [11:0] xfer_stride_bytes; // @[TensorUtil.scala 285:38:@971.4]
  wire [8:0] xfer_stride_pulses; // @[TensorUtil.scala 286:45:@972.4]
  wire  _T_173; // @[TensorUtil.scala 288:21:@973.4]
  wire  _T_175; // @[TensorUtil.scala 289:10:@974.4]
  wire  _T_176; // @[TensorUtil.scala 288:29:@975.4]
  wire [16:0] _T_178; // @[TensorUtil.scala 290:24:@976.4]
  wire [16:0] _T_179; // @[TensorUtil.scala 290:24:@977.4]
  wire [15:0] _T_180; // @[TensorUtil.scala 290:24:@978.4]
  wire  _T_181; // @[TensorUtil.scala 290:10:@979.4]
  wire  stride; // @[TensorUtil.scala 289:18:@980.4]
  wire  _T_184; // @[TensorUtil.scala 292:35:@982.4]
  wire  split; // @[TensorUtil.scala 292:28:@983.4]
  wire [16:0] _GEN_32; // @[TensorUtil.scala 296:16:@986.6]
  wire  _T_185; // @[TensorUtil.scala 296:16:@986.6]
  wire [9:0] _T_188; // @[TensorUtil.scala 300:31:@992.8]
  wire [9:0] _T_189; // @[TensorUtil.scala 300:31:@993.8]
  wire [8:0] _T_190; // @[TensorUtil.scala 300:31:@994.8]
  wire [17:0] _T_191; // @[TensorUtil.scala 301:21:@996.8]
  wire [17:0] _T_192; // @[TensorUtil.scala 301:21:@997.8]
  wire [16:0] _T_193; // @[TensorUtil.scala 301:21:@998.8]
  wire [16:0] _GEN_0; // @[TensorUtil.scala 296:36:@987.6]
  wire [16:0] _GEN_1; // @[TensorUtil.scala 296:36:@987.6]
  wire  _T_194; // @[TensorUtil.scala 303:25:@1003.6]
  wire [16:0] _GEN_34; // @[TensorUtil.scala 305:16:@1006.8]
  wire  _T_195; // @[TensorUtil.scala 305:16:@1006.8]
  wire [9:0] _T_198; // @[TensorUtil.scala 309:33:@1012.10]
  wire [9:0] _T_199; // @[TensorUtil.scala 309:33:@1013.10]
  wire [8:0] _T_200; // @[TensorUtil.scala 309:33:@1014.10]
  wire [17:0] _T_201; // @[TensorUtil.scala 310:21:@1016.10]
  wire [17:0] _T_202; // @[TensorUtil.scala 310:21:@1017.10]
  wire [16:0] _T_203; // @[TensorUtil.scala 310:21:@1018.10]
  wire [16:0] _GEN_2; // @[TensorUtil.scala 305:38:@1007.8]
  wire [16:0] _GEN_3; // @[TensorUtil.scala 305:38:@1007.8]
  wire  _T_204; // @[TensorUtil.scala 312:25:@1023.8]
  wire [15:0] _GEN_36; // @[TensorUtil.scala 314:15:@1026.10]
  wire  _T_205; // @[TensorUtil.scala 314:15:@1026.10]
  wire [9:0] _T_208; // @[TensorUtil.scala 318:32:@1032.12]
  wire [9:0] _T_209; // @[TensorUtil.scala 318:32:@1033.12]
  wire [8:0] _T_210; // @[TensorUtil.scala 318:32:@1034.12]
  wire [16:0] _T_211; // @[TensorUtil.scala 319:20:@1036.12]
  wire [16:0] _T_212; // @[TensorUtil.scala 319:20:@1037.12]
  wire [15:0] _T_213; // @[TensorUtil.scala 319:20:@1038.12]
  wire [15:0] _GEN_4; // @[TensorUtil.scala 314:36:@1027.10]
  wire [15:0] _GEN_5; // @[TensorUtil.scala 314:36:@1027.10]
  wire [31:0] _GEN_6; // @[TensorUtil.scala 312:35:@1024.8]
  wire [15:0] _GEN_7; // @[TensorUtil.scala 312:35:@1024.8]
  wire [15:0] _GEN_8; // @[TensorUtil.scala 312:35:@1024.8]
  wire [31:0] _GEN_9; // @[TensorUtil.scala 303:36:@1004.6]
  wire [16:0] _GEN_10; // @[TensorUtil.scala 303:36:@1004.6]
  wire [16:0] _GEN_11; // @[TensorUtil.scala 303:36:@1004.6]
  wire [16:0] _GEN_13; // @[TensorUtil.scala 294:18:@984.4]
  wire [16:0] _GEN_14; // @[TensorUtil.scala 294:18:@984.4]
  wire [8:0] _T_216; // @[TensorUtil.scala 326:18:@1047.8]
  wire [7:0] _T_217; // @[TensorUtil.scala 326:18:@1048.8]
  wire [7:0] _GEN_15; // @[TensorUtil.scala 325:26:@1046.6]
  wire  _T_219; // @[TensorUtil.scala 331:25:@1055.6]
  wire [16:0] _T_221; // @[TensorUtil.scala 332:18:@1057.8]
  wire [15:0] _T_222; // @[TensorUtil.scala 332:18:@1058.8]
  wire [15:0] _GEN_17; // @[TensorUtil.scala 331:36:@1056.6]
  wire [31:0] _GEN_19; // @[TensorUtil.scala 341:24:@1071.10]
  wire [31:0] _GEN_20; // @[TensorUtil.scala 341:24:@1071.10]
  wire [31:0] _GEN_21; // @[TensorUtil.scala 339:17:@1067.8]
  wire [31:0] _GEN_22; // @[TensorUtil.scala 339:17:@1067.8]
  wire [31:0] _GEN_23; // @[TensorUtil.scala 338:26:@1066.6]
  wire [31:0] _GEN_24; // @[TensorUtil.scala 338:26:@1066.6]
  wire [35:0] _GEN_25; // @[TensorUtil.scala 335:18:@1061.4]
  wire [35:0] _GEN_26; // @[TensorUtil.scala 335:18:@1061.4]
  wire  _T_232; // @[TensorUtil.scala 354:10:@1088.4]
  assign dec_dram_offset = io_inst[56:25]; // @[TensorUtil.scala 251:29:@857.4]
  assign dec_ysize = io_inst[79:64]; // @[TensorUtil.scala 251:29:@861.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 251:29:@863.4]
  assign dec_xstride = io_inst[111:96]; // @[TensorUtil.scala 251:29:@865.4]
  assign _GEN_27 = {{1'd0}, dec_xsize}; // @[TensorUtil.scala 269:26:@944.4]
  assign _T_154 = _GEN_27 << 1; // @[TensorUtil.scala 269:26:@944.4]
  assign _T_156 = _T_154 - 17'h1; // @[TensorUtil.scala 269:51:@945.4]
  assign _T_157 = $unsigned(_T_156); // @[TensorUtil.scala 269:51:@946.4]
  assign xsize = _T_157[16:0]; // @[TensorUtil.scala 269:51:@947.4]
  assign _GEN_28 = {{4'd0}, dec_xstride}; // @[TensorUtil.scala 275:35:@950.4]
  assign xstride_bytes = _GEN_28 << 4; // @[TensorUtil.scala 275:35:@950.4]
  assign _GEN_29 = {{4'd0}, dec_dram_offset}; // @[TensorUtil.scala 277:66:@951.4]
  assign _T_160 = _GEN_29 << 4; // @[TensorUtil.scala 277:66:@951.4]
  assign _T_161 = 36'hffffffff & _T_160; // @[TensorUtil.scala 277:47:@952.4]
  assign _GEN_30 = {{4'd0}, io_baddr}; // @[TensorUtil.scala 277:33:@953.4]
  assign xfer_init_addr = _GEN_30 | _T_161; // @[TensorUtil.scala 277:33:@953.4]
  assign _T_162 = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@954.4]
  assign xfer_split_addr = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@955.4]
  assign _GEN_31 = {{12'd0}, xstride_bytes}; // @[TensorUtil.scala 279:32:@956.4]
  assign _T_163 = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@956.4]
  assign xfer_stride_addr = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@957.4]
  assign _GEN_12 = xfer_init_addr % 36'h800; // @[TensorUtil.scala 281:55:@958.4]
  assign _T_164 = _GEN_12[11:0]; // @[TensorUtil.scala 281:55:@958.4]
  assign _T_165 = 12'h800 - _T_164; // @[TensorUtil.scala 281:38:@959.4]
  assign _T_166 = $unsigned(_T_165); // @[TensorUtil.scala 281:38:@960.4]
  assign xfer_init_bytes = _T_166[11:0]; // @[TensorUtil.scala 281:38:@961.4]
  assign xfer_init_pulses = xfer_init_bytes[11:3]; // @[TensorUtil.scala 282:43:@962.4]
  assign _GEN_16 = xfer_split_addr % 32'h800; // @[TensorUtil.scala 283:56:@963.4]
  assign _T_167 = _GEN_16[11:0]; // @[TensorUtil.scala 283:56:@963.4]
  assign _T_168 = 12'h800 - _T_167; // @[TensorUtil.scala 283:38:@964.4]
  assign _T_169 = $unsigned(_T_168); // @[TensorUtil.scala 283:38:@965.4]
  assign xfer_split_bytes = _T_169[11:0]; // @[TensorUtil.scala 283:38:@966.4]
  assign xfer_split_pulses = xfer_split_bytes[11:3]; // @[TensorUtil.scala 284:44:@967.4]
  assign _GEN_18 = xfer_stride_addr % 32'h800; // @[TensorUtil.scala 285:57:@968.4]
  assign _T_170 = _GEN_18[11:0]; // @[TensorUtil.scala 285:57:@968.4]
  assign _T_171 = 12'h800 - _T_170; // @[TensorUtil.scala 285:38:@969.4]
  assign _T_172 = $unsigned(_T_171); // @[TensorUtil.scala 285:38:@970.4]
  assign xfer_stride_bytes = _T_172[11:0]; // @[TensorUtil.scala 285:38:@971.4]
  assign xfer_stride_pulses = xfer_stride_bytes[11:3]; // @[TensorUtil.scala 286:45:@972.4]
  assign _T_173 = xcnt == len; // @[TensorUtil.scala 288:21:@973.4]
  assign _T_175 = xrem == 16'h0; // @[TensorUtil.scala 289:10:@974.4]
  assign _T_176 = _T_173 & _T_175; // @[TensorUtil.scala 288:29:@975.4]
  assign _T_178 = dec_ysize - 16'h1; // @[TensorUtil.scala 290:24:@976.4]
  assign _T_179 = $unsigned(_T_178); // @[TensorUtil.scala 290:24:@977.4]
  assign _T_180 = _T_179[15:0]; // @[TensorUtil.scala 290:24:@978.4]
  assign _T_181 = ycnt != _T_180; // @[TensorUtil.scala 290:10:@979.4]
  assign stride = _T_176 & _T_181; // @[TensorUtil.scala 289:18:@980.4]
  assign _T_184 = xrem != 16'h0; // @[TensorUtil.scala 292:35:@982.4]
  assign split = _T_173 & _T_184; // @[TensorUtil.scala 292:28:@983.4]
  assign _GEN_32 = {{8'd0}, xfer_init_pulses}; // @[TensorUtil.scala 296:16:@986.6]
  assign _T_185 = xsize < _GEN_32; // @[TensorUtil.scala 296:16:@986.6]
  assign _T_188 = xfer_init_pulses - 9'h1; // @[TensorUtil.scala 300:31:@992.8]
  assign _T_189 = $unsigned(_T_188); // @[TensorUtil.scala 300:31:@993.8]
  assign _T_190 = _T_189[8:0]; // @[TensorUtil.scala 300:31:@994.8]
  assign _T_191 = xsize - _GEN_32; // @[TensorUtil.scala 301:21:@996.8]
  assign _T_192 = $unsigned(_T_191); // @[TensorUtil.scala 301:21:@997.8]
  assign _T_193 = _T_192[16:0]; // @[TensorUtil.scala 301:21:@998.8]
  assign _GEN_0 = _T_185 ? xsize : {{8'd0}, _T_190}; // @[TensorUtil.scala 296:36:@987.6]
  assign _GEN_1 = _T_185 ? 17'h0 : _T_193; // @[TensorUtil.scala 296:36:@987.6]
  assign _T_194 = io_xupdate & stride; // @[TensorUtil.scala 303:25:@1003.6]
  assign _GEN_34 = {{8'd0}, xfer_stride_pulses}; // @[TensorUtil.scala 305:16:@1006.8]
  assign _T_195 = xsize < _GEN_34; // @[TensorUtil.scala 305:16:@1006.8]
  assign _T_198 = xfer_stride_pulses - 9'h1; // @[TensorUtil.scala 309:33:@1012.10]
  assign _T_199 = $unsigned(_T_198); // @[TensorUtil.scala 309:33:@1013.10]
  assign _T_200 = _T_199[8:0]; // @[TensorUtil.scala 309:33:@1014.10]
  assign _T_201 = xsize - _GEN_34; // @[TensorUtil.scala 310:21:@1016.10]
  assign _T_202 = $unsigned(_T_201); // @[TensorUtil.scala 310:21:@1017.10]
  assign _T_203 = _T_202[16:0]; // @[TensorUtil.scala 310:21:@1018.10]
  assign _GEN_2 = _T_195 ? xsize : {{8'd0}, _T_200}; // @[TensorUtil.scala 305:38:@1007.8]
  assign _GEN_3 = _T_195 ? 17'h0 : _T_203; // @[TensorUtil.scala 305:38:@1007.8]
  assign _T_204 = io_xupdate & split; // @[TensorUtil.scala 312:25:@1023.8]
  assign _GEN_36 = {{7'd0}, xfer_split_pulses}; // @[TensorUtil.scala 314:15:@1026.10]
  assign _T_205 = xrem < _GEN_36; // @[TensorUtil.scala 314:15:@1026.10]
  assign _T_208 = xfer_split_pulses - 9'h1; // @[TensorUtil.scala 318:32:@1032.12]
  assign _T_209 = $unsigned(_T_208); // @[TensorUtil.scala 318:32:@1033.12]
  assign _T_210 = _T_209[8:0]; // @[TensorUtil.scala 318:32:@1034.12]
  assign _T_211 = xrem - _GEN_36; // @[TensorUtil.scala 319:20:@1036.12]
  assign _T_212 = $unsigned(_T_211); // @[TensorUtil.scala 319:20:@1037.12]
  assign _T_213 = _T_212[15:0]; // @[TensorUtil.scala 319:20:@1038.12]
  assign _GEN_4 = _T_205 ? xrem : {{7'd0}, _T_210}; // @[TensorUtil.scala 314:36:@1027.10]
  assign _GEN_5 = _T_205 ? 16'h0 : _T_213; // @[TensorUtil.scala 314:36:@1027.10]
  assign _GEN_6 = _T_204 ? {{20'd0}, xfer_split_bytes} : xfer_bytes; // @[TensorUtil.scala 312:35:@1024.8]
  assign _GEN_7 = _T_204 ? _GEN_4 : {{8'd0}, len}; // @[TensorUtil.scala 312:35:@1024.8]
  assign _GEN_8 = _T_204 ? _GEN_5 : xrem; // @[TensorUtil.scala 312:35:@1024.8]
  assign _GEN_9 = _T_194 ? {{20'd0}, xfer_stride_bytes} : _GEN_6; // @[TensorUtil.scala 303:36:@1004.6]
  assign _GEN_10 = _T_194 ? _GEN_2 : {{1'd0}, _GEN_7}; // @[TensorUtil.scala 303:36:@1004.6]
  assign _GEN_11 = _T_194 ? _GEN_3 : {{1'd0}, _GEN_8}; // @[TensorUtil.scala 303:36:@1004.6]
  assign _GEN_13 = io_start ? _GEN_0 : _GEN_10; // @[TensorUtil.scala 294:18:@984.4]
  assign _GEN_14 = io_start ? _GEN_1 : _GEN_11; // @[TensorUtil.scala 294:18:@984.4]
  assign _T_216 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@1047.8]
  assign _T_217 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@1048.8]
  assign _GEN_15 = io_xupdate ? _T_217 : xcnt; // @[TensorUtil.scala 325:26:@1046.6]
  assign _T_219 = io_yupdate & stride; // @[TensorUtil.scala 331:25:@1055.6]
  assign _T_221 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@1057.8]
  assign _T_222 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@1058.8]
  assign _GEN_17 = _T_219 ? _T_222 : ycnt; // @[TensorUtil.scala 331:36:@1056.6]
  assign _GEN_19 = stride ? xfer_stride_addr : caddr; // @[TensorUtil.scala 341:24:@1071.10]
  assign _GEN_20 = stride ? xfer_stride_addr : baddr; // @[TensorUtil.scala 341:24:@1071.10]
  assign _GEN_21 = split ? xfer_split_addr : _GEN_19; // @[TensorUtil.scala 339:17:@1067.8]
  assign _GEN_22 = split ? baddr : _GEN_20; // @[TensorUtil.scala 339:17:@1067.8]
  assign _GEN_23 = io_yupdate ? _GEN_21 : caddr; // @[TensorUtil.scala 338:26:@1066.6]
  assign _GEN_24 = io_yupdate ? _GEN_22 : baddr; // @[TensorUtil.scala 338:26:@1066.6]
  assign _GEN_25 = io_start ? xfer_init_addr : {{4'd0}, _GEN_23}; // @[TensorUtil.scala 335:18:@1061.4]
  assign _GEN_26 = io_start ? xfer_init_addr : {{4'd0}, _GEN_24}; // @[TensorUtil.scala 335:18:@1061.4]
  assign _T_232 = ycnt == _T_180; // @[TensorUtil.scala 354:10:@1088.4]
  assign io_done = _T_176 & _T_232; // @[TensorUtil.scala 352:11:@1090.4]
  assign io_stride = _T_176 & _T_181; // @[TensorUtil.scala 347:13:@1076.4]
  assign io_split = _T_173 & _T_184; // @[TensorUtil.scala 348:12:@1077.4]
  assign io_addr = caddr; // @[TensorUtil.scala 350:11:@1080.4]
  assign io_len = len; // @[TensorUtil.scala 351:10:@1081.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  caddr = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  baddr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  len = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  xcnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xrem = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ycnt = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  xfer_bytes = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    caddr <= _GEN_25[31:0];
    baddr <= _GEN_26[31:0];
    len <= _GEN_13[7:0];
    if (io_xinit) begin
      xcnt <= 8'h0;
    end else begin
      if (io_xupdate) begin
        xcnt <= _T_217;
      end
    end
    xrem <= _GEN_14[15:0];
    if (io_start) begin
      ycnt <= 16'h0;
    end else begin
      if (_T_219) begin
        ycnt <= _T_222;
      end
    end
    if (io_start) begin
      xfer_bytes <= {{20'd0}, xfer_init_bytes};
    end else begin
      if (_T_194) begin
        xfer_bytes <= {{20'd0}, xfer_stride_bytes};
      end else begin
        if (_T_204) begin
          xfer_bytes <= {{20'd0}, xfer_split_bytes};
        end
      end
    end
  end
endmodule
module TensorPadCtrl( // @[:@1092.2]
  input          clock, // @[:@1093.4]
  input          reset, // @[:@1094.4]
  input          io_start, // @[:@1095.4]
  output         io_done, // @[:@1095.4]
  input  [127:0] io_inst // @[:@1095.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@1120.4]
  wire [3:0] dec_ypad_0; // @[TensorUtil.scala 173:29:@1124.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@1128.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@1130.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@1132.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@1133.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@1134.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@1135.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@1136.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@1136.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@1137.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@1138.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@1138.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@1139.4]
  wire [16:0] _GEN_12; // @[TensorUtil.scala 182:46:@1140.4]
  wire [16:0] _T_39; // @[TensorUtil.scala 182:46:@1140.4]
  wire [17:0] _T_41; // @[TensorUtil.scala 182:71:@1141.4]
  wire [17:0] _T_42; // @[TensorUtil.scala 182:71:@1142.4]
  wire [16:0] xval; // @[TensorUtil.scala 182:71:@1143.4]
  wire  _T_44; // @[TensorUtil.scala 190:22:@1144.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 190:42:@1145.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 190:42:@1146.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 190:42:@1147.4]
  wire [3:0] yval; // @[TensorUtil.scala 190:10:@1148.4]
  reg  state; // @[TensorUtil.scala 197:22:@1149.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@1150.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@1152.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@1159.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@1160.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@1161.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@1162.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@1158.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@1151.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@1166.4]
  wire [16:0] _GEN_4; // @[TensorUtil.scala 212:25:@1167.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@1173.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@1180.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@1181.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@1179.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@1185.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@1186.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@1193.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@1195.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@1196.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@1194.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@1201.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@1120.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorUtil.scala 173:29:@1124.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@1128.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@1130.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@1136.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@1136.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@1137.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@1138.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@1138.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@1139.4]
  assign _GEN_12 = {{1'd0}, _T_38}; // @[TensorUtil.scala 182:46:@1140.4]
  assign _T_39 = _GEN_12 << 1; // @[TensorUtil.scala 182:46:@1140.4]
  assign _T_41 = _T_39 - 17'h1; // @[TensorUtil.scala 182:71:@1141.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@1142.4]
  assign xval = _T_42[16:0]; // @[TensorUtil.scala 182:71:@1143.4]
  assign _T_44 = dec_ypad_0 != 4'h0; // @[TensorUtil.scala 190:22:@1144.4]
  assign _T_46 = dec_ypad_0 - 4'h1; // @[TensorUtil.scala 190:42:@1145.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 190:42:@1146.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 190:42:@1147.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 190:10:@1148.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@1150.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@1152.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@1159.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@1160.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@1161.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@1162.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@1158.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@1151.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@1166.4]
  assign _GEN_4 = _T_56 ? xval : {{1'd0}, xmax}; // @[TensorUtil.scala 212:25:@1167.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@1173.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1180.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1181.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@1179.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@1185.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@1186.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@1193.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@1195.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@1196.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@1194.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@1201.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@1204.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_1( // @[:@1206.2]
  input          clock, // @[:@1207.4]
  input          reset, // @[:@1208.4]
  input          io_start, // @[:@1209.4]
  output         io_done, // @[:@1209.4]
  input  [127:0] io_inst // @[:@1209.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@1234.4]
  wire [3:0] dec_ypad_1; // @[TensorUtil.scala 173:29:@1240.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@1242.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@1244.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@1246.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@1247.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@1248.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@1249.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@1250.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@1250.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@1251.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@1252.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@1252.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@1253.4]
  wire [16:0] _GEN_12; // @[TensorUtil.scala 182:46:@1254.4]
  wire [16:0] _T_39; // @[TensorUtil.scala 182:46:@1254.4]
  wire [17:0] _T_41; // @[TensorUtil.scala 182:71:@1255.4]
  wire [17:0] _T_42; // @[TensorUtil.scala 182:71:@1256.4]
  wire [16:0] xval; // @[TensorUtil.scala 182:71:@1257.4]
  wire  _T_44; // @[TensorUtil.scala 192:22:@1258.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 192:42:@1259.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 192:42:@1260.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 192:42:@1261.4]
  wire [3:0] yval; // @[TensorUtil.scala 192:10:@1262.4]
  reg  state; // @[TensorUtil.scala 197:22:@1263.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@1264.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@1266.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@1273.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@1274.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@1275.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@1276.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@1272.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@1265.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@1280.4]
  wire [16:0] _GEN_4; // @[TensorUtil.scala 212:25:@1281.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@1287.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@1294.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@1295.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@1293.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@1299.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@1300.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@1307.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@1309.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@1310.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@1308.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@1315.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@1234.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorUtil.scala 173:29:@1240.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@1242.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@1244.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@1250.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@1250.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@1251.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@1252.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@1252.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@1253.4]
  assign _GEN_12 = {{1'd0}, _T_38}; // @[TensorUtil.scala 182:46:@1254.4]
  assign _T_39 = _GEN_12 << 1; // @[TensorUtil.scala 182:46:@1254.4]
  assign _T_41 = _T_39 - 17'h1; // @[TensorUtil.scala 182:71:@1255.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@1256.4]
  assign xval = _T_42[16:0]; // @[TensorUtil.scala 182:71:@1257.4]
  assign _T_44 = dec_ypad_1 != 4'h0; // @[TensorUtil.scala 192:22:@1258.4]
  assign _T_46 = dec_ypad_1 - 4'h1; // @[TensorUtil.scala 192:42:@1259.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 192:42:@1260.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 192:42:@1261.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 192:10:@1262.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@1264.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@1266.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@1273.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@1274.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@1275.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@1276.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@1272.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@1265.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@1280.4]
  assign _GEN_4 = _T_56 ? xval : {{1'd0}, xmax}; // @[TensorUtil.scala 212:25:@1281.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@1287.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1294.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1295.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@1293.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@1299.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@1300.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@1307.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@1309.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@1310.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@1308.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@1315.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@1318.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_2( // @[:@1320.2]
  input          clock, // @[:@1321.4]
  input          reset, // @[:@1322.4]
  input          io_start, // @[:@1323.4]
  output         io_done, // @[:@1323.4]
  input  [127:0] io_inst // @[:@1323.4]
);
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@1356.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@1360.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@1362.4]
  reg [31:0] _RAND_1;
  wire [4:0] _GEN_10; // @[TensorUtil.scala 184:19:@1364.4]
  wire [4:0] _T_35; // @[TensorUtil.scala 184:19:@1364.4]
  wire [5:0] _T_37; // @[TensorUtil.scala 184:44:@1365.4]
  wire [5:0] _T_38; // @[TensorUtil.scala 184:44:@1366.4]
  wire [4:0] xval; // @[TensorUtil.scala 184:44:@1367.4]
  reg  state; // @[TensorUtil.scala 197:22:@1368.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@1369.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@1371.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@1379.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@1381.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@1377.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@1370.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@1385.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@1392.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@1399.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@1400.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@1398.6]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@1356.4]
  assign _GEN_10 = {{1'd0}, dec_xpad_0}; // @[TensorUtil.scala 184:19:@1364.4]
  assign _T_35 = _GEN_10 << 1; // @[TensorUtil.scala 184:19:@1364.4]
  assign _T_37 = _T_35 - 5'h1; // @[TensorUtil.scala 184:44:@1365.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 184:44:@1366.4]
  assign xval = _T_38[4:0]; // @[TensorUtil.scala 184:44:@1367.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@1369.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@1371.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@1379.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@1381.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@1377.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@1370.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@1385.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@1392.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1399.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1400.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@1398.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@1423.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{11'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_3( // @[:@1425.2]
  input          clock, // @[:@1426.4]
  input          reset, // @[:@1427.4]
  input          io_start, // @[:@1428.4]
  output         io_done, // @[:@1428.4]
  input  [127:0] io_inst // @[:@1428.4]
);
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@1463.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@1465.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@1467.4]
  reg [31:0] _RAND_1;
  wire [4:0] _GEN_10; // @[TensorUtil.scala 186:19:@1469.4]
  wire [4:0] _T_35; // @[TensorUtil.scala 186:19:@1469.4]
  wire [5:0] _T_37; // @[TensorUtil.scala 186:44:@1470.4]
  wire [5:0] _T_38; // @[TensorUtil.scala 186:44:@1471.4]
  wire [4:0] xval; // @[TensorUtil.scala 186:44:@1472.4]
  reg  state; // @[TensorUtil.scala 197:22:@1473.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@1474.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@1476.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@1484.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@1486.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@1482.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@1475.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@1490.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@1497.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@1504.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@1505.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@1503.6]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@1463.4]
  assign _GEN_10 = {{1'd0}, dec_xpad_1}; // @[TensorUtil.scala 186:19:@1469.4]
  assign _T_35 = _GEN_10 << 1; // @[TensorUtil.scala 186:19:@1469.4]
  assign _T_37 = _T_35 - 5'h1; // @[TensorUtil.scala 186:44:@1470.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 186:44:@1471.4]
  assign xval = _T_38[4:0]; // @[TensorUtil.scala 186:44:@1472.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@1474.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@1476.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@1484.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@1486.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@1482.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@1475.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@1490.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@1497.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1504.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1505.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@1503.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@1528.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{11'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorLoad( // @[:@1530.2]
  input          clock, // @[:@1531.4]
  input          reset, // @[:@1532.4]
  input          io_start, // @[:@1533.4]
  output         io_done, // @[:@1533.4]
  input  [127:0] io_inst, // @[:@1533.4]
  input  [31:0]  io_baddr, // @[:@1533.4]
  input          io_vme_rd_cmd_ready, // @[:@1533.4]
  output         io_vme_rd_cmd_valid, // @[:@1533.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@1533.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@1533.4]
  output         io_vme_rd_data_ready, // @[:@1533.4]
  input          io_vme_rd_data_valid, // @[:@1533.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@1533.4]
  input          io_tensor_rd_idx_valid, // @[:@1533.4]
  input  [10:0]  io_tensor_rd_idx_bits, // @[:@1533.4]
  output         io_tensor_rd_data_valid, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_0, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_1, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_2, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_3, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_4, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_5, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_6, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_7, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_8, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_9, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_10, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_11, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_12, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_13, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_14, // @[:@1533.4]
  output [7:0]   io_tensor_rd_data_bits_0_15 // @[:@1533.4]
);
  wire  dataCtrl_clock; // @[TensorLoad.scala 52:24:@1570.4]
  wire  dataCtrl_io_start; // @[TensorLoad.scala 52:24:@1570.4]
  wire  dataCtrl_io_done; // @[TensorLoad.scala 52:24:@1570.4]
  wire [127:0] dataCtrl_io_inst; // @[TensorLoad.scala 52:24:@1570.4]
  wire [31:0] dataCtrl_io_baddr; // @[TensorLoad.scala 52:24:@1570.4]
  wire  dataCtrl_io_xinit; // @[TensorLoad.scala 52:24:@1570.4]
  wire  dataCtrl_io_xupdate; // @[TensorLoad.scala 52:24:@1570.4]
  wire  dataCtrl_io_yupdate; // @[TensorLoad.scala 52:24:@1570.4]
  wire  dataCtrl_io_stride; // @[TensorLoad.scala 52:24:@1570.4]
  wire  dataCtrl_io_split; // @[TensorLoad.scala 52:24:@1570.4]
  wire [31:0] dataCtrl_io_addr; // @[TensorLoad.scala 52:24:@1570.4]
  wire [7:0] dataCtrl_io_len; // @[TensorLoad.scala 52:24:@1570.4]
  wire  yPadCtrl0_clock; // @[TensorLoad.scala 55:25:@1574.4]
  wire  yPadCtrl0_reset; // @[TensorLoad.scala 55:25:@1574.4]
  wire  yPadCtrl0_io_start; // @[TensorLoad.scala 55:25:@1574.4]
  wire  yPadCtrl0_io_done; // @[TensorLoad.scala 55:25:@1574.4]
  wire [127:0] yPadCtrl0_io_inst; // @[TensorLoad.scala 55:25:@1574.4]
  wire  yPadCtrl1_clock; // @[TensorLoad.scala 56:25:@1577.4]
  wire  yPadCtrl1_reset; // @[TensorLoad.scala 56:25:@1577.4]
  wire  yPadCtrl1_io_start; // @[TensorLoad.scala 56:25:@1577.4]
  wire  yPadCtrl1_io_done; // @[TensorLoad.scala 56:25:@1577.4]
  wire [127:0] yPadCtrl1_io_inst; // @[TensorLoad.scala 56:25:@1577.4]
  wire  xPadCtrl0_clock; // @[TensorLoad.scala 57:25:@1580.4]
  wire  xPadCtrl0_reset; // @[TensorLoad.scala 57:25:@1580.4]
  wire  xPadCtrl0_io_start; // @[TensorLoad.scala 57:25:@1580.4]
  wire  xPadCtrl0_io_done; // @[TensorLoad.scala 57:25:@1580.4]
  wire [127:0] xPadCtrl0_io_inst; // @[TensorLoad.scala 57:25:@1580.4]
  wire  xPadCtrl1_clock; // @[TensorLoad.scala 58:25:@1583.4]
  wire  xPadCtrl1_reset; // @[TensorLoad.scala 58:25:@1583.4]
  wire  xPadCtrl1_io_start; // @[TensorLoad.scala 58:25:@1583.4]
  wire  xPadCtrl1_io_done; // @[TensorLoad.scala 58:25:@1583.4]
  wire [127:0] xPadCtrl1_io_inst; // @[TensorLoad.scala 58:25:@1583.4]
  reg [63:0] tensorFile_0_0 [0:2047]; // @[TensorLoad.scala 222:16:@1853.4]
  reg [63:0] _RAND_0;
  wire [63:0] tensorFile_0_0_rdata_0_data; // @[TensorLoad.scala 222:16:@1853.4]
  wire [10:0] tensorFile_0_0_rdata_0_addr; // @[TensorLoad.scala 222:16:@1853.4]
  wire [63:0] tensorFile_0_0__T_866_data; // @[TensorLoad.scala 222:16:@1853.4]
  wire [10:0] tensorFile_0_0__T_866_addr; // @[TensorLoad.scala 222:16:@1853.4]
  wire  tensorFile_0_0__T_866_mask; // @[TensorLoad.scala 222:16:@1853.4]
  wire  tensorFile_0_0__T_866_en; // @[TensorLoad.scala 222:16:@1853.4]
  reg [63:0] tensorFile_0_1 [0:2047]; // @[TensorLoad.scala 222:16:@1853.4]
  reg [63:0] _RAND_1;
  wire [63:0] tensorFile_0_1_rdata_0_data; // @[TensorLoad.scala 222:16:@1853.4]
  wire [10:0] tensorFile_0_1_rdata_0_addr; // @[TensorLoad.scala 222:16:@1853.4]
  wire [63:0] tensorFile_0_1__T_866_data; // @[TensorLoad.scala 222:16:@1853.4]
  wire [10:0] tensorFile_0_1__T_866_addr; // @[TensorLoad.scala 222:16:@1853.4]
  wire  tensorFile_0_1__T_866_mask; // @[TensorLoad.scala 222:16:@1853.4]
  wire  tensorFile_0_1__T_866_en; // @[TensorLoad.scala 222:16:@1853.4]
  wire [15:0] dec_sram_offset; // @[TensorLoad.scala 51:29:@1550.4]
  wire [15:0] dec_xsize; // @[TensorLoad.scala 51:29:@1558.4]
  wire [3:0] dec_ypad_0; // @[TensorLoad.scala 51:29:@1562.4]
  wire [3:0] dec_ypad_1; // @[TensorLoad.scala 51:29:@1564.4]
  wire [3:0] dec_xpad_0; // @[TensorLoad.scala 51:29:@1566.4]
  wire [3:0] dec_xpad_1; // @[TensorLoad.scala 51:29:@1568.4]
  reg  dataCtrlDone; // @[TensorLoad.scala 54:29:@1573.4]
  reg [31:0] _RAND_2;
  reg  tag; // @[TensorLoad.scala 60:16:@1586.4]
  reg [31:0] _RAND_3;
  reg [2:0] state; // @[TensorLoad.scala 65:22:@1588.4]
  reg [31:0] _RAND_4;
  wire  _T_614; // @[Conditional.scala 37:30:@1589.4]
  wire  _T_616; // @[TensorLoad.scala 71:25:@1592.8]
  wire  _T_618; // @[TensorLoad.scala 73:31:@1597.10]
  wire [2:0] _GEN_0; // @[TensorLoad.scala 73:40:@1598.10]
  wire [2:0] _GEN_1; // @[TensorLoad.scala 71:34:@1593.8]
  wire [2:0] _GEN_2; // @[TensorLoad.scala 70:22:@1591.6]
  wire  _T_619; // @[Conditional.scala 37:30:@1607.6]
  wire [2:0] _GEN_4; // @[TensorLoad.scala 81:31:@1609.8]
  wire  _T_622; // @[Conditional.scala 37:30:@1620.8]
  wire [2:0] _GEN_5; // @[TensorLoad.scala 90:31:@1622.10]
  wire  _T_623; // @[Conditional.scala 37:30:@1627.10]
  wire [2:0] _GEN_6; // @[TensorLoad.scala 95:33:@1629.12]
  wire  _T_624; // @[Conditional.scala 37:30:@1634.12]
  wire  _T_626; // @[TensorLoad.scala 102:27:@1638.18]
  wire  _T_628; // @[TensorLoad.scala 104:33:@1643.20]
  wire [2:0] _GEN_7; // @[TensorLoad.scala 104:42:@1644.20]
  wire [2:0] _GEN_8; // @[TensorLoad.scala 102:36:@1639.18]
  wire [2:0] _GEN_10; // @[TensorLoad.scala 110:36:@1654.20]
  wire [2:0] _GEN_11; // @[TensorLoad.scala 117:39:@1667.20]
  wire [2:0] _GEN_12; // @[TensorLoad.scala 109:40:@1652.18]
  wire [2:0] _GEN_13; // @[TensorLoad.scala 101:32:@1637.16]
  wire [2:0] _GEN_14; // @[TensorLoad.scala 100:34:@1636.14]
  wire  _T_633; // @[Conditional.scala 37:30:@1673.14]
  wire [2:0] _GEN_17; // @[TensorLoad.scala 124:28:@1676.18]
  wire [2:0] _GEN_18; // @[TensorLoad.scala 123:31:@1675.16]
  wire  _T_638; // @[Conditional.scala 37:30:@1697.16]
  wire  _T_639; // @[TensorLoad.scala 140:30:@1699.18]
  wire [2:0] _GEN_19; // @[TensorLoad.scala 140:47:@1700.18]
  wire [2:0] _GEN_20; // @[Conditional.scala 39:67:@1698.16]
  wire [2:0] _GEN_21; // @[Conditional.scala 39:67:@1674.14]
  wire [2:0] _GEN_22; // @[Conditional.scala 39:67:@1635.12]
  wire [2:0] _GEN_23; // @[Conditional.scala 39:67:@1628.10]
  wire [2:0] _GEN_24; // @[Conditional.scala 39:67:@1621.8]
  wire [2:0] _GEN_25; // @[Conditional.scala 39:67:@1608.6]
  wire [2:0] _GEN_26; // @[Conditional.scala 40:58:@1590.4]
  wire  _T_640; // @[TensorLoad.scala 147:30:@1704.4]
  wire  _T_641; // @[TensorLoad.scala 147:40:@1705.4]
  wire  _T_643; // @[Decoupled.scala 37:37:@1711.4]
  wire  _T_648; // @[TensorLoad.scala 156:36:@1721.6]
  wire  _GEN_27; // @[TensorLoad.scala 156:57:@1722.6]
  wire  _GEN_28; // @[TensorLoad.scala 154:25:@1716.4]
  wire  _T_653; // @[TensorLoad.scala 161:44:@1727.4]
  wire  _T_660; // @[TensorLoad.scala 164:61:@1733.4]
  wire  _T_661; // @[TensorLoad.scala 164:48:@1734.4]
  wire  _T_662; // @[TensorLoad.scala 165:14:@1735.4]
  wire  _T_663; // @[TensorLoad.scala 165:25:@1736.4]
  wire  _T_664; // @[TensorLoad.scala 165:45:@1737.4]
  wire  _T_665; // @[TensorLoad.scala 164:70:@1738.4]
  wire  _T_671; // @[TensorLoad.scala 169:14:@1744.4]
  wire  _T_672; // @[TensorLoad.scala 169:25:@1745.4]
  wire  _T_673; // @[TensorLoad.scala 168:35:@1746.4]
  wire  _T_675; // @[TensorLoad.scala 170:32:@1748.4]
  wire  _T_676; // @[TensorLoad.scala 170:30:@1749.4]
  wire  _T_677; // @[TensorLoad.scala 170:46:@1750.4]
  wire  _T_680; // @[TensorLoad.scala 170:67:@1752.4]
  wire  _T_681; // @[TensorLoad.scala 169:46:@1753.4]
  wire  _T_685; // @[TensorLoad.scala 171:45:@1757.4]
  wire  _T_686; // @[TensorLoad.scala 170:89:@1758.4]
  wire  _T_691; // @[TensorLoad.scala 173:44:@1763.4]
  wire  _T_692; // @[TensorLoad.scala 174:28:@1764.4]
  wire  _T_693; // @[TensorLoad.scala 174:46:@1765.4]
  wire  _T_696; // @[TensorLoad.scala 174:67:@1767.4]
  wire  _T_697; // @[TensorLoad.scala 174:25:@1768.4]
  wire  _T_699; // @[TensorLoad.scala 182:32:@1775.4]
  wire  _T_702; // @[TensorLoad.scala 190:11:@1782.4]
  wire  _T_703; // @[TensorLoad.scala 189:36:@1783.4]
  wire  _T_705; // @[TensorLoad.scala 190:22:@1785.4]
  wire  _T_706; // @[TensorLoad.scala 192:11:@1786.4]
  wire  isZeroPad; // @[TensorLoad.scala 191:22:@1787.4]
  wire  _T_709; // @[TensorLoad.scala 194:24:@1790.4]
  wire  _T_712; // @[TensorLoad.scala 194:46:@1792.4]
  wire  _T_715; // @[TensorLoad.scala 196:36:@1798.6]
  wire [1:0] _T_717; // @[TensorLoad.scala 197:16:@1800.8]
  wire  _T_718; // @[TensorLoad.scala 197:16:@1801.8]
  wire  _GEN_29; // @[TensorLoad.scala 196:50:@1799.6]
  wire  _T_732; // @[TensorLoad.scala 202:51:@1817.6]
  reg [10:0] waddr_cur; // @[TensorLoad.scala 206:22:@1823.4]
  reg [31:0] _RAND_5;
  reg [10:0] waddr_nxt; // @[TensorLoad.scala 207:22:@1824.4]
  reg [31:0] _RAND_6;
  wire [11:0] _T_748; // @[TensorLoad.scala 215:28:@1838.8]
  wire [10:0] _T_749; // @[TensorLoad.scala 215:28:@1839.8]
  wire  _T_751; // @[TensorLoad.scala 216:33:@1844.8]
  wire [15:0] _GEN_66; // @[TensorLoad.scala 217:28:@1846.10]
  wire [16:0] _T_752; // @[TensorLoad.scala 217:28:@1846.10]
  wire [15:0] _T_753; // @[TensorLoad.scala 217:28:@1847.10]
  wire [15:0] _GEN_33; // @[TensorLoad.scala 216:59:@1845.8]
  wire [15:0] _GEN_34; // @[TensorLoad.scala 216:59:@1845.8]
  wire [15:0] _GEN_35; // @[TensorLoad.scala 214:3:@1837.6]
  wire [15:0] _GEN_36; // @[TensorLoad.scala 214:3:@1837.6]
  wire [15:0] _GEN_37; // @[TensorLoad.scala 208:25:@1826.4]
  wire [15:0] _GEN_38; // @[TensorLoad.scala 208:25:@1826.4]
  wire  wmask_0_0; // @[TensorLoad.scala 235:26:@1859.4]
  wire [63:0] wdata_0_0; // @[TensorLoad.scala 236:25:@1861.4]
  reg  rvalid; // @[TensorLoad.scala 252:23:@1910.4]
  reg [31:0] _RAND_7;
  wire  _GEN_51; // @[TensorLoad.scala 256:26:@1915.4]
  wire [127:0] _T_887; // @[TensorLoad.scala 259:38:@1921.4]
  wire  _T_1035; // @[TensorLoad.scala 263:96:@1977.4]
  wire  done_no_pad; // @[TensorLoad.scala 263:83:@1978.4]
  wire  done_x_pad; // @[TensorLoad.scala 264:72:@1983.4]
  wire  _T_1042; // @[TensorLoad.scala 265:37:@1985.4]
  wire  done_y_pad; // @[TensorLoad.scala 265:52:@1986.4]
  wire  _T_1043; // @[TensorLoad.scala 266:26:@1987.4]
  reg [10:0] tensorFile_0_0_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [10:0] tensorFile_0_1_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_9;
  TensorDataCtrl dataCtrl ( // @[TensorLoad.scala 52:24:@1570.4]
    .clock(dataCtrl_clock),
    .io_start(dataCtrl_io_start),
    .io_done(dataCtrl_io_done),
    .io_inst(dataCtrl_io_inst),
    .io_baddr(dataCtrl_io_baddr),
    .io_xinit(dataCtrl_io_xinit),
    .io_xupdate(dataCtrl_io_xupdate),
    .io_yupdate(dataCtrl_io_yupdate),
    .io_stride(dataCtrl_io_stride),
    .io_split(dataCtrl_io_split),
    .io_addr(dataCtrl_io_addr),
    .io_len(dataCtrl_io_len)
  );
  TensorPadCtrl yPadCtrl0 ( // @[TensorLoad.scala 55:25:@1574.4]
    .clock(yPadCtrl0_clock),
    .reset(yPadCtrl0_reset),
    .io_start(yPadCtrl0_io_start),
    .io_done(yPadCtrl0_io_done),
    .io_inst(yPadCtrl0_io_inst)
  );
  TensorPadCtrl_1 yPadCtrl1 ( // @[TensorLoad.scala 56:25:@1577.4]
    .clock(yPadCtrl1_clock),
    .reset(yPadCtrl1_reset),
    .io_start(yPadCtrl1_io_start),
    .io_done(yPadCtrl1_io_done),
    .io_inst(yPadCtrl1_io_inst)
  );
  TensorPadCtrl_2 xPadCtrl0 ( // @[TensorLoad.scala 57:25:@1580.4]
    .clock(xPadCtrl0_clock),
    .reset(xPadCtrl0_reset),
    .io_start(xPadCtrl0_io_start),
    .io_done(xPadCtrl0_io_done),
    .io_inst(xPadCtrl0_io_inst)
  );
  TensorPadCtrl_3 xPadCtrl1 ( // @[TensorLoad.scala 58:25:@1583.4]
    .clock(xPadCtrl1_clock),
    .reset(xPadCtrl1_reset),
    .io_start(xPadCtrl1_io_start),
    .io_done(xPadCtrl1_io_done),
    .io_inst(xPadCtrl1_io_inst)
  );
  assign tensorFile_0_0_rdata_0_addr = tensorFile_0_0_rdata_0_addr_pipe_0;
  assign tensorFile_0_0_rdata_0_data = tensorFile_0_0[tensorFile_0_0_rdata_0_addr]; // @[TensorLoad.scala 222:16:@1853.4]
  assign tensorFile_0_0__T_866_data = _T_640 ? 64'h0 : wdata_0_0;
  assign tensorFile_0_0__T_866_addr = _T_640 ? 11'h0 : waddr_cur;
  assign tensorFile_0_0__T_866_mask = _T_640 ? 1'h1 : wmask_0_0;
  assign tensorFile_0_0__T_866_en = _T_640 ? 1'h0 : _T_715;
  assign tensorFile_0_1_rdata_0_addr = tensorFile_0_1_rdata_0_addr_pipe_0;
  assign tensorFile_0_1_rdata_0_data = tensorFile_0_1[tensorFile_0_1_rdata_0_addr]; // @[TensorLoad.scala 222:16:@1853.4]
  assign tensorFile_0_1__T_866_data = _T_640 ? 64'h0 : wdata_0_0;
  assign tensorFile_0_1__T_866_addr = _T_640 ? 11'h0 : waddr_cur;
  assign tensorFile_0_1__T_866_mask = _T_640 ? 1'h1 : tag;
  assign tensorFile_0_1__T_866_en = _T_640 ? 1'h0 : _T_715;
  assign dec_sram_offset = io_inst[24:9]; // @[TensorLoad.scala 51:29:@1550.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorLoad.scala 51:29:@1558.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorLoad.scala 51:29:@1562.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorLoad.scala 51:29:@1564.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorLoad.scala 51:29:@1566.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorLoad.scala 51:29:@1568.4]
  assign _T_614 = 3'h0 == state; // @[Conditional.scala 37:30:@1589.4]
  assign _T_616 = dec_ypad_0 != 4'h0; // @[TensorLoad.scala 71:25:@1592.8]
  assign _T_618 = dec_xpad_0 != 4'h0; // @[TensorLoad.scala 73:31:@1597.10]
  assign _GEN_0 = _T_618 ? 3'h2 : 3'h3; // @[TensorLoad.scala 73:40:@1598.10]
  assign _GEN_1 = _T_616 ? 3'h1 : _GEN_0; // @[TensorLoad.scala 71:34:@1593.8]
  assign _GEN_2 = io_start ? _GEN_1 : state; // @[TensorLoad.scala 70:22:@1591.6]
  assign _T_619 = 3'h1 == state; // @[Conditional.scala 37:30:@1607.6]
  assign _GEN_4 = yPadCtrl0_io_done ? _GEN_0 : state; // @[TensorLoad.scala 81:31:@1609.8]
  assign _T_622 = 3'h2 == state; // @[Conditional.scala 37:30:@1620.8]
  assign _GEN_5 = xPadCtrl0_io_done ? 3'h3 : state; // @[TensorLoad.scala 90:31:@1622.10]
  assign _T_623 = 3'h3 == state; // @[Conditional.scala 37:30:@1627.10]
  assign _GEN_6 = io_vme_rd_cmd_ready ? 3'h4 : state; // @[TensorLoad.scala 95:33:@1629.12]
  assign _T_624 = 3'h4 == state; // @[Conditional.scala 37:30:@1634.12]
  assign _T_626 = dec_xpad_1 != 4'h0; // @[TensorLoad.scala 102:27:@1638.18]
  assign _T_628 = dec_ypad_1 != 4'h0; // @[TensorLoad.scala 104:33:@1643.20]
  assign _GEN_7 = _T_628 ? 3'h6 : 3'h0; // @[TensorLoad.scala 104:42:@1644.20]
  assign _GEN_8 = _T_626 ? 3'h5 : _GEN_7; // @[TensorLoad.scala 102:36:@1639.18]
  assign _GEN_10 = _T_626 ? 3'h5 : _GEN_0; // @[TensorLoad.scala 110:36:@1654.20]
  assign _GEN_11 = dataCtrl_io_split ? 3'h3 : state; // @[TensorLoad.scala 117:39:@1667.20]
  assign _GEN_12 = dataCtrl_io_stride ? _GEN_10 : _GEN_11; // @[TensorLoad.scala 109:40:@1652.18]
  assign _GEN_13 = dataCtrl_io_done ? _GEN_8 : _GEN_12; // @[TensorLoad.scala 101:32:@1637.16]
  assign _GEN_14 = io_vme_rd_data_valid ? _GEN_13 : state; // @[TensorLoad.scala 100:34:@1636.14]
  assign _T_633 = 3'h5 == state; // @[Conditional.scala 37:30:@1673.14]
  assign _GEN_17 = dataCtrlDone ? _GEN_7 : _GEN_0; // @[TensorLoad.scala 124:28:@1676.18]
  assign _GEN_18 = xPadCtrl1_io_done ? _GEN_17 : state; // @[TensorLoad.scala 123:31:@1675.16]
  assign _T_638 = 3'h6 == state; // @[Conditional.scala 37:30:@1697.16]
  assign _T_639 = yPadCtrl1_io_done & dataCtrlDone; // @[TensorLoad.scala 140:30:@1699.18]
  assign _GEN_19 = _T_639 ? 3'h0 : state; // @[TensorLoad.scala 140:47:@1700.18]
  assign _GEN_20 = _T_638 ? _GEN_19 : state; // @[Conditional.scala 39:67:@1698.16]
  assign _GEN_21 = _T_633 ? _GEN_18 : _GEN_20; // @[Conditional.scala 39:67:@1674.14]
  assign _GEN_22 = _T_624 ? _GEN_14 : _GEN_21; // @[Conditional.scala 39:67:@1635.12]
  assign _GEN_23 = _T_623 ? _GEN_6 : _GEN_22; // @[Conditional.scala 39:67:@1628.10]
  assign _GEN_24 = _T_622 ? _GEN_5 : _GEN_23; // @[Conditional.scala 39:67:@1621.8]
  assign _GEN_25 = _T_619 ? _GEN_4 : _GEN_24; // @[Conditional.scala 39:67:@1608.6]
  assign _GEN_26 = _T_614 ? _GEN_2 : _GEN_25; // @[Conditional.scala 40:58:@1590.4]
  assign _T_640 = state == 3'h0; // @[TensorLoad.scala 147:30:@1704.4]
  assign _T_641 = _T_640 & io_start; // @[TensorLoad.scala 147:40:@1705.4]
  assign _T_643 = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[Decoupled.scala 37:37:@1711.4]
  assign _T_648 = _T_643 & dataCtrl_io_done; // @[TensorLoad.scala 156:36:@1721.6]
  assign _GEN_27 = _T_648 ? 1'h1 : dataCtrlDone; // @[TensorLoad.scala 156:57:@1722.6]
  assign _GEN_28 = _T_640 ? 1'h0 : _GEN_27; // @[TensorLoad.scala 154:25:@1716.4]
  assign _T_653 = _T_616 & _T_640; // @[TensorLoad.scala 161:44:@1727.4]
  assign _T_660 = dec_xpad_1 == 4'h0; // @[TensorLoad.scala 164:61:@1733.4]
  assign _T_661 = _T_648 & _T_660; // @[TensorLoad.scala 164:48:@1734.4]
  assign _T_662 = state == 3'h5; // @[TensorLoad.scala 165:14:@1735.4]
  assign _T_663 = _T_662 & xPadCtrl1_io_done; // @[TensorLoad.scala 165:25:@1736.4]
  assign _T_664 = _T_663 & dataCtrlDone; // @[TensorLoad.scala 165:45:@1737.4]
  assign _T_665 = _T_661 | _T_664; // @[TensorLoad.scala 164:70:@1738.4]
  assign _T_671 = state == 3'h1; // @[TensorLoad.scala 169:14:@1744.4]
  assign _T_672 = _T_671 & yPadCtrl0_io_done; // @[TensorLoad.scala 169:25:@1745.4]
  assign _T_673 = _T_641 | _T_672; // @[TensorLoad.scala 168:35:@1746.4]
  assign _T_675 = ~ dataCtrlDone; // @[TensorLoad.scala 170:32:@1748.4]
  assign _T_676 = _T_643 & _T_675; // @[TensorLoad.scala 170:30:@1749.4]
  assign _T_677 = _T_676 & dataCtrl_io_stride; // @[TensorLoad.scala 170:46:@1750.4]
  assign _T_680 = _T_677 & _T_660; // @[TensorLoad.scala 170:67:@1752.4]
  assign _T_681 = _T_673 | _T_680; // @[TensorLoad.scala 169:46:@1753.4]
  assign _T_685 = _T_663 & _T_675; // @[TensorLoad.scala 171:45:@1757.4]
  assign _T_686 = _T_681 | _T_685; // @[TensorLoad.scala 170:89:@1758.4]
  assign _T_691 = _T_626 & _T_643; // @[TensorLoad.scala 173:44:@1763.4]
  assign _T_692 = ~ dataCtrl_io_done; // @[TensorLoad.scala 174:28:@1764.4]
  assign _T_693 = _T_692 & dataCtrl_io_stride; // @[TensorLoad.scala 174:46:@1765.4]
  assign _T_696 = _T_693 & _T_626; // @[TensorLoad.scala 174:67:@1767.4]
  assign _T_697 = dataCtrl_io_done | _T_696; // @[TensorLoad.scala 174:25:@1768.4]
  assign _T_699 = state == 3'h3; // @[TensorLoad.scala 182:32:@1775.4]
  assign _T_702 = state == 3'h2; // @[TensorLoad.scala 190:11:@1782.4]
  assign _T_703 = _T_671 | _T_702; // @[TensorLoad.scala 189:36:@1783.4]
  assign _T_705 = _T_703 | _T_662; // @[TensorLoad.scala 190:22:@1785.4]
  assign _T_706 = state == 3'h6; // @[TensorLoad.scala 192:11:@1786.4]
  assign isZeroPad = _T_705 | _T_706; // @[TensorLoad.scala 191:22:@1787.4]
  assign _T_709 = _T_640 | _T_699; // @[TensorLoad.scala 194:24:@1790.4]
  assign _T_712 = _T_709 | tag; // @[TensorLoad.scala 194:46:@1792.4]
  assign _T_715 = _T_643 | isZeroPad; // @[TensorLoad.scala 196:36:@1798.6]
  assign _T_717 = tag + 1'h1; // @[TensorLoad.scala 197:16:@1800.8]
  assign _T_718 = tag + 1'h1; // @[TensorLoad.scala 197:16:@1801.8]
  assign _GEN_29 = _T_715 ? _T_718 : tag; // @[TensorLoad.scala 196:50:@1799.6]
  assign _T_732 = _T_715 & tag; // @[TensorLoad.scala 202:51:@1817.6]
  assign _T_748 = waddr_cur + 11'h1; // @[TensorLoad.scala 215:28:@1838.8]
  assign _T_749 = waddr_cur + 11'h1; // @[TensorLoad.scala 215:28:@1839.8]
  assign _T_751 = dataCtrl_io_stride & _T_643; // @[TensorLoad.scala 216:33:@1844.8]
  assign _GEN_66 = {{5'd0}, waddr_nxt}; // @[TensorLoad.scala 217:28:@1846.10]
  assign _T_752 = _GEN_66 + dec_xsize; // @[TensorLoad.scala 217:28:@1846.10]
  assign _T_753 = _GEN_66 + dec_xsize; // @[TensorLoad.scala 217:28:@1847.10]
  assign _GEN_33 = _T_751 ? _T_753 : {{5'd0}, waddr_cur}; // @[TensorLoad.scala 216:59:@1845.8]
  assign _GEN_34 = _T_751 ? _T_753 : {{5'd0}, waddr_nxt}; // @[TensorLoad.scala 216:59:@1845.8]
  assign _GEN_35 = _T_732 ? {{5'd0}, _T_749} : _GEN_33; // @[TensorLoad.scala 214:3:@1837.6]
  assign _GEN_36 = _T_732 ? {{5'd0}, waddr_nxt} : _GEN_34; // @[TensorLoad.scala 214:3:@1837.6]
  assign _GEN_37 = _T_640 ? dec_sram_offset : _GEN_35; // @[TensorLoad.scala 208:25:@1826.4]
  assign _GEN_38 = _T_640 ? dec_sram_offset : _GEN_36; // @[TensorLoad.scala 208:25:@1826.4]
  assign wmask_0_0 = tag == 1'h0; // @[TensorLoad.scala 235:26:@1859.4]
  assign wdata_0_0 = isZeroPad ? 64'h0 : io_vme_rd_data_bits; // @[TensorLoad.scala 236:25:@1861.4]
  assign _GEN_51 = io_tensor_rd_idx_valid; // @[TensorLoad.scala 256:26:@1915.4]
  assign _T_887 = {tensorFile_0_1_rdata_0_data,tensorFile_0_0_rdata_0_data}; // @[TensorLoad.scala 259:38:@1921.4]
  assign _T_1035 = dec_ypad_1 == 4'h0; // @[TensorLoad.scala 263:96:@1977.4]
  assign done_no_pad = _T_661 & _T_1035; // @[TensorLoad.scala 263:83:@1978.4]
  assign done_x_pad = _T_664 & _T_1035; // @[TensorLoad.scala 264:72:@1983.4]
  assign _T_1042 = _T_706 & dataCtrlDone; // @[TensorLoad.scala 265:37:@1985.4]
  assign done_y_pad = _T_1042 & yPadCtrl1_io_done; // @[TensorLoad.scala 265:52:@1986.4]
  assign _T_1043 = done_no_pad | done_x_pad; // @[TensorLoad.scala 266:26:@1987.4]
  assign io_done = _T_1043 | done_y_pad; // @[TensorLoad.scala 266:11:@1989.4]
  assign io_vme_rd_cmd_valid = state == 3'h3; // @[TensorLoad.scala 182:23:@1776.4]
  assign io_vme_rd_cmd_bits_addr = dataCtrl_io_addr; // @[TensorLoad.scala 183:27:@1777.4]
  assign io_vme_rd_cmd_bits_len = dataCtrl_io_len; // @[TensorLoad.scala 184:26:@1778.4]
  assign io_vme_rd_data_ready = state == 3'h4; // @[TensorLoad.scala 186:24:@1780.4]
  assign io_tensor_rd_data_valid = rvalid; // @[TensorLoad.scala 253:27:@1912.4]
  assign io_tensor_rd_data_bits_0_0 = _T_887[7:0]; // @[TensorLoad.scala 259:33:@1957.4]
  assign io_tensor_rd_data_bits_0_1 = _T_887[15:8]; // @[TensorLoad.scala 259:33:@1958.4]
  assign io_tensor_rd_data_bits_0_2 = _T_887[23:16]; // @[TensorLoad.scala 259:33:@1959.4]
  assign io_tensor_rd_data_bits_0_3 = _T_887[31:24]; // @[TensorLoad.scala 259:33:@1960.4]
  assign io_tensor_rd_data_bits_0_4 = _T_887[39:32]; // @[TensorLoad.scala 259:33:@1961.4]
  assign io_tensor_rd_data_bits_0_5 = _T_887[47:40]; // @[TensorLoad.scala 259:33:@1962.4]
  assign io_tensor_rd_data_bits_0_6 = _T_887[55:48]; // @[TensorLoad.scala 259:33:@1963.4]
  assign io_tensor_rd_data_bits_0_7 = _T_887[63:56]; // @[TensorLoad.scala 259:33:@1964.4]
  assign io_tensor_rd_data_bits_0_8 = _T_887[71:64]; // @[TensorLoad.scala 259:33:@1965.4]
  assign io_tensor_rd_data_bits_0_9 = _T_887[79:72]; // @[TensorLoad.scala 259:33:@1966.4]
  assign io_tensor_rd_data_bits_0_10 = _T_887[87:80]; // @[TensorLoad.scala 259:33:@1967.4]
  assign io_tensor_rd_data_bits_0_11 = _T_887[95:88]; // @[TensorLoad.scala 259:33:@1968.4]
  assign io_tensor_rd_data_bits_0_12 = _T_887[103:96]; // @[TensorLoad.scala 259:33:@1969.4]
  assign io_tensor_rd_data_bits_0_13 = _T_887[111:104]; // @[TensorLoad.scala 259:33:@1970.4]
  assign io_tensor_rd_data_bits_0_14 = _T_887[119:112]; // @[TensorLoad.scala 259:33:@1971.4]
  assign io_tensor_rd_data_bits_0_15 = _T_887[127:120]; // @[TensorLoad.scala 259:33:@1972.4]
  assign dataCtrl_clock = clock; // @[:@1571.4]
  assign dataCtrl_io_start = _T_640 & io_start; // @[TensorLoad.scala 147:21:@1706.4]
  assign dataCtrl_io_inst = io_inst; // @[TensorLoad.scala 148:20:@1707.4]
  assign dataCtrl_io_baddr = io_baddr; // @[TensorLoad.scala 149:21:@1708.4]
  assign dataCtrl_io_xinit = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[TensorLoad.scala 150:21:@1710.4]
  assign dataCtrl_io_xupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 151:23:@1712.4]
  assign dataCtrl_io_yupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 152:23:@1714.4]
  assign yPadCtrl0_clock = clock; // @[:@1575.4]
  assign yPadCtrl0_reset = reset; // @[:@1576.4]
  assign yPadCtrl0_io_start = _T_653 & io_start; // @[TensorLoad.scala 161:22:@1729.4]
  assign yPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 176:21:@1771.4]
  assign yPadCtrl1_clock = clock; // @[:@1578.4]
  assign yPadCtrl1_reset = reset; // @[:@1579.4]
  assign yPadCtrl1_io_start = _T_628 & _T_665; // @[TensorLoad.scala 163:22:@1740.4]
  assign yPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 177:21:@1772.4]
  assign xPadCtrl0_clock = clock; // @[:@1581.4]
  assign xPadCtrl0_reset = reset; // @[:@1582.4]
  assign xPadCtrl0_io_start = _T_618 & _T_686; // @[TensorLoad.scala 167:22:@1760.4]
  assign xPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 178:21:@1773.4]
  assign xPadCtrl1_clock = clock; // @[:@1584.4]
  assign xPadCtrl1_reset = reset; // @[:@1585.4]
  assign xPadCtrl1_io_start = _T_691 & _T_697; // @[TensorLoad.scala 173:22:@1770.4]
  assign xPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 179:21:@1774.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_0[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_1[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  dataCtrlDone = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  tag = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  waddr_cur = _RAND_5[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  waddr_nxt = _RAND_6[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rvalid = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tensorFile_0_0_rdata_0_addr_pipe_0 = _RAND_8[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  tensorFile_0_1_rdata_0_addr_pipe_0 = _RAND_9[10:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tensorFile_0_0__T_866_en & tensorFile_0_0__T_866_mask) begin
      tensorFile_0_0[tensorFile_0_0__T_866_addr] <= tensorFile_0_0__T_866_data; // @[TensorLoad.scala 222:16:@1853.4]
    end
    if(tensorFile_0_1__T_866_en & tensorFile_0_1__T_866_mask) begin
      tensorFile_0_1[tensorFile_0_1__T_866_addr] <= tensorFile_0_1__T_866_data; // @[TensorLoad.scala 222:16:@1853.4]
    end
    if (reset) begin
      dataCtrlDone <= 1'h0;
    end else begin
      if (_T_640) begin
        dataCtrlDone <= 1'h0;
      end else begin
        if (_T_648) begin
          dataCtrlDone <= 1'h1;
        end
      end
    end
    if (_T_712) begin
      tag <= 1'h0;
    end else begin
      if (_T_715) begin
        tag <= _T_718;
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_614) begin
        if (io_start) begin
          if (_T_616) begin
            state <= 3'h1;
          end else begin
            if (_T_618) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end
      end else begin
        if (_T_619) begin
          if (yPadCtrl0_io_done) begin
            if (_T_618) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end else begin
          if (_T_622) begin
            if (xPadCtrl0_io_done) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_623) begin
              if (io_vme_rd_cmd_ready) begin
                state <= 3'h4;
              end
            end else begin
              if (_T_624) begin
                if (io_vme_rd_data_valid) begin
                  if (dataCtrl_io_done) begin
                    if (_T_626) begin
                      state <= 3'h5;
                    end else begin
                      if (_T_628) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end
                  end else begin
                    if (dataCtrl_io_stride) begin
                      if (_T_626) begin
                        state <= 3'h5;
                      end else begin
                        if (_T_618) begin
                          state <= 3'h2;
                        end else begin
                          state <= 3'h3;
                        end
                      end
                    end else begin
                      if (dataCtrl_io_split) begin
                        state <= 3'h3;
                      end
                    end
                  end
                end
              end else begin
                if (_T_633) begin
                  if (xPadCtrl1_io_done) begin
                    if (dataCtrlDone) begin
                      if (_T_628) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end else begin
                      if (_T_618) begin
                        state <= 3'h2;
                      end else begin
                        state <= 3'h3;
                      end
                    end
                  end
                end else begin
                  if (_T_638) begin
                    if (_T_639) begin
                      state <= 3'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    waddr_cur <= _GEN_37[10:0];
    waddr_nxt <= _GEN_38[10:0];
    rvalid <= io_tensor_rd_idx_valid;
    if (_GEN_51) begin
      tensorFile_0_0_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_51) begin
      tensorFile_0_1_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
  end
endmodule
module TensorDataCtrl_1( // @[:@1991.2]
  input          clock, // @[:@1992.4]
  input          io_start, // @[:@1994.4]
  output         io_done, // @[:@1994.4]
  input  [127:0] io_inst, // @[:@1994.4]
  input  [31:0]  io_baddr, // @[:@1994.4]
  input          io_xinit, // @[:@1994.4]
  input          io_xupdate, // @[:@1994.4]
  input          io_yupdate, // @[:@1994.4]
  output         io_stride, // @[:@1994.4]
  output         io_split, // @[:@1994.4]
  output [31:0]  io_addr, // @[:@1994.4]
  output [7:0]   io_len // @[:@1994.4]
);
  wire [31:0] dec_dram_offset; // @[TensorUtil.scala 251:29:@2013.4]
  wire [15:0] dec_ysize; // @[TensorUtil.scala 251:29:@2017.4]
  wire [15:0] dec_xsize; // @[TensorUtil.scala 251:29:@2019.4]
  wire [15:0] dec_xstride; // @[TensorUtil.scala 251:29:@2021.4]
  reg [31:0] caddr; // @[TensorUtil.scala 253:18:@2031.4]
  reg [31:0] _RAND_0;
  reg [31:0] baddr; // @[TensorUtil.scala 254:18:@2032.4]
  reg [31:0] _RAND_1;
  reg [7:0] len; // @[TensorUtil.scala 255:16:@2033.4]
  reg [31:0] _RAND_2;
  reg [7:0] xcnt; // @[TensorUtil.scala 267:17:@2098.4]
  reg [31:0] _RAND_3;
  reg [15:0] xrem; // @[TensorUtil.scala 268:17:@2099.4]
  reg [31:0] _RAND_4;
  wire [20:0] _GEN_27; // @[TensorUtil.scala 269:26:@2100.4]
  wire [20:0] _T_154; // @[TensorUtil.scala 269:26:@2100.4]
  wire [21:0] _T_156; // @[TensorUtil.scala 269:51:@2101.4]
  wire [21:0] _T_157; // @[TensorUtil.scala 269:51:@2102.4]
  wire [20:0] xsize; // @[TensorUtil.scala 269:51:@2103.4]
  reg [15:0] ycnt; // @[TensorUtil.scala 271:17:@2104.4]
  reg [31:0] _RAND_5;
  reg [31:0] xfer_bytes; // @[TensorUtil.scala 273:23:@2105.4]
  reg [31:0] _RAND_6;
  wire [23:0] _GEN_28; // @[TensorUtil.scala 275:35:@2106.4]
  wire [23:0] xstride_bytes; // @[TensorUtil.scala 275:35:@2106.4]
  wire [39:0] _GEN_29; // @[TensorUtil.scala 277:66:@2107.4]
  wire [39:0] _T_160; // @[TensorUtil.scala 277:66:@2107.4]
  wire [39:0] _T_161; // @[TensorUtil.scala 277:47:@2108.4]
  wire [39:0] _GEN_30; // @[TensorUtil.scala 277:33:@2109.4]
  wire [39:0] xfer_init_addr; // @[TensorUtil.scala 277:33:@2109.4]
  wire [32:0] _T_162; // @[TensorUtil.scala 278:31:@2110.4]
  wire [31:0] xfer_split_addr; // @[TensorUtil.scala 278:31:@2111.4]
  wire [31:0] _GEN_31; // @[TensorUtil.scala 279:32:@2112.4]
  wire [32:0] _T_163; // @[TensorUtil.scala 279:32:@2112.4]
  wire [31:0] xfer_stride_addr; // @[TensorUtil.scala 279:32:@2113.4]
  wire [39:0] _GEN_12; // @[TensorUtil.scala 281:55:@2114.4]
  wire [11:0] _T_164; // @[TensorUtil.scala 281:55:@2114.4]
  wire [12:0] _T_165; // @[TensorUtil.scala 281:38:@2115.4]
  wire [12:0] _T_166; // @[TensorUtil.scala 281:38:@2116.4]
  wire [11:0] xfer_init_bytes; // @[TensorUtil.scala 281:38:@2117.4]
  wire [8:0] xfer_init_pulses; // @[TensorUtil.scala 282:43:@2118.4]
  wire [31:0] _GEN_16; // @[TensorUtil.scala 283:56:@2119.4]
  wire [11:0] _T_167; // @[TensorUtil.scala 283:56:@2119.4]
  wire [12:0] _T_168; // @[TensorUtil.scala 283:38:@2120.4]
  wire [12:0] _T_169; // @[TensorUtil.scala 283:38:@2121.4]
  wire [11:0] xfer_split_bytes; // @[TensorUtil.scala 283:38:@2122.4]
  wire [8:0] xfer_split_pulses; // @[TensorUtil.scala 284:44:@2123.4]
  wire [31:0] _GEN_18; // @[TensorUtil.scala 285:57:@2124.4]
  wire [11:0] _T_170; // @[TensorUtil.scala 285:57:@2124.4]
  wire [12:0] _T_171; // @[TensorUtil.scala 285:38:@2125.4]
  wire [12:0] _T_172; // @[TensorUtil.scala 285:38:@2126.4]
  wire [11:0] xfer_stride_bytes; // @[TensorUtil.scala 285:38:@2127.4]
  wire [8:0] xfer_stride_pulses; // @[TensorUtil.scala 286:45:@2128.4]
  wire  _T_173; // @[TensorUtil.scala 288:21:@2129.4]
  wire  _T_175; // @[TensorUtil.scala 289:10:@2130.4]
  wire  _T_176; // @[TensorUtil.scala 288:29:@2131.4]
  wire [16:0] _T_178; // @[TensorUtil.scala 290:24:@2132.4]
  wire [16:0] _T_179; // @[TensorUtil.scala 290:24:@2133.4]
  wire [15:0] _T_180; // @[TensorUtil.scala 290:24:@2134.4]
  wire  _T_181; // @[TensorUtil.scala 290:10:@2135.4]
  wire  stride; // @[TensorUtil.scala 289:18:@2136.4]
  wire  _T_184; // @[TensorUtil.scala 292:35:@2138.4]
  wire  split; // @[TensorUtil.scala 292:28:@2139.4]
  wire [20:0] _GEN_32; // @[TensorUtil.scala 296:16:@2142.6]
  wire  _T_185; // @[TensorUtil.scala 296:16:@2142.6]
  wire [9:0] _T_188; // @[TensorUtil.scala 300:31:@2148.8]
  wire [9:0] _T_189; // @[TensorUtil.scala 300:31:@2149.8]
  wire [8:0] _T_190; // @[TensorUtil.scala 300:31:@2150.8]
  wire [21:0] _T_191; // @[TensorUtil.scala 301:21:@2152.8]
  wire [21:0] _T_192; // @[TensorUtil.scala 301:21:@2153.8]
  wire [20:0] _T_193; // @[TensorUtil.scala 301:21:@2154.8]
  wire [20:0] _GEN_0; // @[TensorUtil.scala 296:36:@2143.6]
  wire [20:0] _GEN_1; // @[TensorUtil.scala 296:36:@2143.6]
  wire  _T_194; // @[TensorUtil.scala 303:25:@2159.6]
  wire [20:0] _GEN_34; // @[TensorUtil.scala 305:16:@2162.8]
  wire  _T_195; // @[TensorUtil.scala 305:16:@2162.8]
  wire [9:0] _T_198; // @[TensorUtil.scala 309:33:@2168.10]
  wire [9:0] _T_199; // @[TensorUtil.scala 309:33:@2169.10]
  wire [8:0] _T_200; // @[TensorUtil.scala 309:33:@2170.10]
  wire [21:0] _T_201; // @[TensorUtil.scala 310:21:@2172.10]
  wire [21:0] _T_202; // @[TensorUtil.scala 310:21:@2173.10]
  wire [20:0] _T_203; // @[TensorUtil.scala 310:21:@2174.10]
  wire [20:0] _GEN_2; // @[TensorUtil.scala 305:38:@2163.8]
  wire [20:0] _GEN_3; // @[TensorUtil.scala 305:38:@2163.8]
  wire  _T_204; // @[TensorUtil.scala 312:25:@2179.8]
  wire [15:0] _GEN_36; // @[TensorUtil.scala 314:15:@2182.10]
  wire  _T_205; // @[TensorUtil.scala 314:15:@2182.10]
  wire [9:0] _T_208; // @[TensorUtil.scala 318:32:@2188.12]
  wire [9:0] _T_209; // @[TensorUtil.scala 318:32:@2189.12]
  wire [8:0] _T_210; // @[TensorUtil.scala 318:32:@2190.12]
  wire [16:0] _T_211; // @[TensorUtil.scala 319:20:@2192.12]
  wire [16:0] _T_212; // @[TensorUtil.scala 319:20:@2193.12]
  wire [15:0] _T_213; // @[TensorUtil.scala 319:20:@2194.12]
  wire [15:0] _GEN_4; // @[TensorUtil.scala 314:36:@2183.10]
  wire [15:0] _GEN_5; // @[TensorUtil.scala 314:36:@2183.10]
  wire [31:0] _GEN_6; // @[TensorUtil.scala 312:35:@2180.8]
  wire [15:0] _GEN_7; // @[TensorUtil.scala 312:35:@2180.8]
  wire [15:0] _GEN_8; // @[TensorUtil.scala 312:35:@2180.8]
  wire [31:0] _GEN_9; // @[TensorUtil.scala 303:36:@2160.6]
  wire [20:0] _GEN_10; // @[TensorUtil.scala 303:36:@2160.6]
  wire [20:0] _GEN_11; // @[TensorUtil.scala 303:36:@2160.6]
  wire [20:0] _GEN_13; // @[TensorUtil.scala 294:18:@2140.4]
  wire [20:0] _GEN_14; // @[TensorUtil.scala 294:18:@2140.4]
  wire [8:0] _T_216; // @[TensorUtil.scala 326:18:@2203.8]
  wire [7:0] _T_217; // @[TensorUtil.scala 326:18:@2204.8]
  wire [7:0] _GEN_15; // @[TensorUtil.scala 325:26:@2202.6]
  wire  _T_219; // @[TensorUtil.scala 331:25:@2211.6]
  wire [16:0] _T_221; // @[TensorUtil.scala 332:18:@2213.8]
  wire [15:0] _T_222; // @[TensorUtil.scala 332:18:@2214.8]
  wire [15:0] _GEN_17; // @[TensorUtil.scala 331:36:@2212.6]
  wire [31:0] _GEN_19; // @[TensorUtil.scala 341:24:@2227.10]
  wire [31:0] _GEN_20; // @[TensorUtil.scala 341:24:@2227.10]
  wire [31:0] _GEN_21; // @[TensorUtil.scala 339:17:@2223.8]
  wire [31:0] _GEN_22; // @[TensorUtil.scala 339:17:@2223.8]
  wire [31:0] _GEN_23; // @[TensorUtil.scala 338:26:@2222.6]
  wire [31:0] _GEN_24; // @[TensorUtil.scala 338:26:@2222.6]
  wire [39:0] _GEN_25; // @[TensorUtil.scala 335:18:@2217.4]
  wire [39:0] _GEN_26; // @[TensorUtil.scala 335:18:@2217.4]
  wire  _T_232; // @[TensorUtil.scala 354:10:@2244.4]
  assign dec_dram_offset = io_inst[56:25]; // @[TensorUtil.scala 251:29:@2013.4]
  assign dec_ysize = io_inst[79:64]; // @[TensorUtil.scala 251:29:@2017.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 251:29:@2019.4]
  assign dec_xstride = io_inst[111:96]; // @[TensorUtil.scala 251:29:@2021.4]
  assign _GEN_27 = {{5'd0}, dec_xsize}; // @[TensorUtil.scala 269:26:@2100.4]
  assign _T_154 = _GEN_27 << 5; // @[TensorUtil.scala 269:26:@2100.4]
  assign _T_156 = _T_154 - 21'h1; // @[TensorUtil.scala 269:51:@2101.4]
  assign _T_157 = $unsigned(_T_156); // @[TensorUtil.scala 269:51:@2102.4]
  assign xsize = _T_157[20:0]; // @[TensorUtil.scala 269:51:@2103.4]
  assign _GEN_28 = {{8'd0}, dec_xstride}; // @[TensorUtil.scala 275:35:@2106.4]
  assign xstride_bytes = _GEN_28 << 8; // @[TensorUtil.scala 275:35:@2106.4]
  assign _GEN_29 = {{8'd0}, dec_dram_offset}; // @[TensorUtil.scala 277:66:@2107.4]
  assign _T_160 = _GEN_29 << 8; // @[TensorUtil.scala 277:66:@2107.4]
  assign _T_161 = 40'hffffffff & _T_160; // @[TensorUtil.scala 277:47:@2108.4]
  assign _GEN_30 = {{8'd0}, io_baddr}; // @[TensorUtil.scala 277:33:@2109.4]
  assign xfer_init_addr = _GEN_30 | _T_161; // @[TensorUtil.scala 277:33:@2109.4]
  assign _T_162 = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@2110.4]
  assign xfer_split_addr = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@2111.4]
  assign _GEN_31 = {{8'd0}, xstride_bytes}; // @[TensorUtil.scala 279:32:@2112.4]
  assign _T_163 = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@2112.4]
  assign xfer_stride_addr = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@2113.4]
  assign _GEN_12 = xfer_init_addr % 40'h800; // @[TensorUtil.scala 281:55:@2114.4]
  assign _T_164 = _GEN_12[11:0]; // @[TensorUtil.scala 281:55:@2114.4]
  assign _T_165 = 12'h800 - _T_164; // @[TensorUtil.scala 281:38:@2115.4]
  assign _T_166 = $unsigned(_T_165); // @[TensorUtil.scala 281:38:@2116.4]
  assign xfer_init_bytes = _T_166[11:0]; // @[TensorUtil.scala 281:38:@2117.4]
  assign xfer_init_pulses = xfer_init_bytes[11:3]; // @[TensorUtil.scala 282:43:@2118.4]
  assign _GEN_16 = xfer_split_addr % 32'h800; // @[TensorUtil.scala 283:56:@2119.4]
  assign _T_167 = _GEN_16[11:0]; // @[TensorUtil.scala 283:56:@2119.4]
  assign _T_168 = 12'h800 - _T_167; // @[TensorUtil.scala 283:38:@2120.4]
  assign _T_169 = $unsigned(_T_168); // @[TensorUtil.scala 283:38:@2121.4]
  assign xfer_split_bytes = _T_169[11:0]; // @[TensorUtil.scala 283:38:@2122.4]
  assign xfer_split_pulses = xfer_split_bytes[11:3]; // @[TensorUtil.scala 284:44:@2123.4]
  assign _GEN_18 = xfer_stride_addr % 32'h800; // @[TensorUtil.scala 285:57:@2124.4]
  assign _T_170 = _GEN_18[11:0]; // @[TensorUtil.scala 285:57:@2124.4]
  assign _T_171 = 12'h800 - _T_170; // @[TensorUtil.scala 285:38:@2125.4]
  assign _T_172 = $unsigned(_T_171); // @[TensorUtil.scala 285:38:@2126.4]
  assign xfer_stride_bytes = _T_172[11:0]; // @[TensorUtil.scala 285:38:@2127.4]
  assign xfer_stride_pulses = xfer_stride_bytes[11:3]; // @[TensorUtil.scala 286:45:@2128.4]
  assign _T_173 = xcnt == len; // @[TensorUtil.scala 288:21:@2129.4]
  assign _T_175 = xrem == 16'h0; // @[TensorUtil.scala 289:10:@2130.4]
  assign _T_176 = _T_173 & _T_175; // @[TensorUtil.scala 288:29:@2131.4]
  assign _T_178 = dec_ysize - 16'h1; // @[TensorUtil.scala 290:24:@2132.4]
  assign _T_179 = $unsigned(_T_178); // @[TensorUtil.scala 290:24:@2133.4]
  assign _T_180 = _T_179[15:0]; // @[TensorUtil.scala 290:24:@2134.4]
  assign _T_181 = ycnt != _T_180; // @[TensorUtil.scala 290:10:@2135.4]
  assign stride = _T_176 & _T_181; // @[TensorUtil.scala 289:18:@2136.4]
  assign _T_184 = xrem != 16'h0; // @[TensorUtil.scala 292:35:@2138.4]
  assign split = _T_173 & _T_184; // @[TensorUtil.scala 292:28:@2139.4]
  assign _GEN_32 = {{12'd0}, xfer_init_pulses}; // @[TensorUtil.scala 296:16:@2142.6]
  assign _T_185 = xsize < _GEN_32; // @[TensorUtil.scala 296:16:@2142.6]
  assign _T_188 = xfer_init_pulses - 9'h1; // @[TensorUtil.scala 300:31:@2148.8]
  assign _T_189 = $unsigned(_T_188); // @[TensorUtil.scala 300:31:@2149.8]
  assign _T_190 = _T_189[8:0]; // @[TensorUtil.scala 300:31:@2150.8]
  assign _T_191 = xsize - _GEN_32; // @[TensorUtil.scala 301:21:@2152.8]
  assign _T_192 = $unsigned(_T_191); // @[TensorUtil.scala 301:21:@2153.8]
  assign _T_193 = _T_192[20:0]; // @[TensorUtil.scala 301:21:@2154.8]
  assign _GEN_0 = _T_185 ? xsize : {{12'd0}, _T_190}; // @[TensorUtil.scala 296:36:@2143.6]
  assign _GEN_1 = _T_185 ? 21'h0 : _T_193; // @[TensorUtil.scala 296:36:@2143.6]
  assign _T_194 = io_xupdate & stride; // @[TensorUtil.scala 303:25:@2159.6]
  assign _GEN_34 = {{12'd0}, xfer_stride_pulses}; // @[TensorUtil.scala 305:16:@2162.8]
  assign _T_195 = xsize < _GEN_34; // @[TensorUtil.scala 305:16:@2162.8]
  assign _T_198 = xfer_stride_pulses - 9'h1; // @[TensorUtil.scala 309:33:@2168.10]
  assign _T_199 = $unsigned(_T_198); // @[TensorUtil.scala 309:33:@2169.10]
  assign _T_200 = _T_199[8:0]; // @[TensorUtil.scala 309:33:@2170.10]
  assign _T_201 = xsize - _GEN_34; // @[TensorUtil.scala 310:21:@2172.10]
  assign _T_202 = $unsigned(_T_201); // @[TensorUtil.scala 310:21:@2173.10]
  assign _T_203 = _T_202[20:0]; // @[TensorUtil.scala 310:21:@2174.10]
  assign _GEN_2 = _T_195 ? xsize : {{12'd0}, _T_200}; // @[TensorUtil.scala 305:38:@2163.8]
  assign _GEN_3 = _T_195 ? 21'h0 : _T_203; // @[TensorUtil.scala 305:38:@2163.8]
  assign _T_204 = io_xupdate & split; // @[TensorUtil.scala 312:25:@2179.8]
  assign _GEN_36 = {{7'd0}, xfer_split_pulses}; // @[TensorUtil.scala 314:15:@2182.10]
  assign _T_205 = xrem < _GEN_36; // @[TensorUtil.scala 314:15:@2182.10]
  assign _T_208 = xfer_split_pulses - 9'h1; // @[TensorUtil.scala 318:32:@2188.12]
  assign _T_209 = $unsigned(_T_208); // @[TensorUtil.scala 318:32:@2189.12]
  assign _T_210 = _T_209[8:0]; // @[TensorUtil.scala 318:32:@2190.12]
  assign _T_211 = xrem - _GEN_36; // @[TensorUtil.scala 319:20:@2192.12]
  assign _T_212 = $unsigned(_T_211); // @[TensorUtil.scala 319:20:@2193.12]
  assign _T_213 = _T_212[15:0]; // @[TensorUtil.scala 319:20:@2194.12]
  assign _GEN_4 = _T_205 ? xrem : {{7'd0}, _T_210}; // @[TensorUtil.scala 314:36:@2183.10]
  assign _GEN_5 = _T_205 ? 16'h0 : _T_213; // @[TensorUtil.scala 314:36:@2183.10]
  assign _GEN_6 = _T_204 ? {{20'd0}, xfer_split_bytes} : xfer_bytes; // @[TensorUtil.scala 312:35:@2180.8]
  assign _GEN_7 = _T_204 ? _GEN_4 : {{8'd0}, len}; // @[TensorUtil.scala 312:35:@2180.8]
  assign _GEN_8 = _T_204 ? _GEN_5 : xrem; // @[TensorUtil.scala 312:35:@2180.8]
  assign _GEN_9 = _T_194 ? {{20'd0}, xfer_stride_bytes} : _GEN_6; // @[TensorUtil.scala 303:36:@2160.6]
  assign _GEN_10 = _T_194 ? _GEN_2 : {{5'd0}, _GEN_7}; // @[TensorUtil.scala 303:36:@2160.6]
  assign _GEN_11 = _T_194 ? _GEN_3 : {{5'd0}, _GEN_8}; // @[TensorUtil.scala 303:36:@2160.6]
  assign _GEN_13 = io_start ? _GEN_0 : _GEN_10; // @[TensorUtil.scala 294:18:@2140.4]
  assign _GEN_14 = io_start ? _GEN_1 : _GEN_11; // @[TensorUtil.scala 294:18:@2140.4]
  assign _T_216 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@2203.8]
  assign _T_217 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@2204.8]
  assign _GEN_15 = io_xupdate ? _T_217 : xcnt; // @[TensorUtil.scala 325:26:@2202.6]
  assign _T_219 = io_yupdate & stride; // @[TensorUtil.scala 331:25:@2211.6]
  assign _T_221 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@2213.8]
  assign _T_222 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@2214.8]
  assign _GEN_17 = _T_219 ? _T_222 : ycnt; // @[TensorUtil.scala 331:36:@2212.6]
  assign _GEN_19 = stride ? xfer_stride_addr : caddr; // @[TensorUtil.scala 341:24:@2227.10]
  assign _GEN_20 = stride ? xfer_stride_addr : baddr; // @[TensorUtil.scala 341:24:@2227.10]
  assign _GEN_21 = split ? xfer_split_addr : _GEN_19; // @[TensorUtil.scala 339:17:@2223.8]
  assign _GEN_22 = split ? baddr : _GEN_20; // @[TensorUtil.scala 339:17:@2223.8]
  assign _GEN_23 = io_yupdate ? _GEN_21 : caddr; // @[TensorUtil.scala 338:26:@2222.6]
  assign _GEN_24 = io_yupdate ? _GEN_22 : baddr; // @[TensorUtil.scala 338:26:@2222.6]
  assign _GEN_25 = io_start ? xfer_init_addr : {{8'd0}, _GEN_23}; // @[TensorUtil.scala 335:18:@2217.4]
  assign _GEN_26 = io_start ? xfer_init_addr : {{8'd0}, _GEN_24}; // @[TensorUtil.scala 335:18:@2217.4]
  assign _T_232 = ycnt == _T_180; // @[TensorUtil.scala 354:10:@2244.4]
  assign io_done = _T_176 & _T_232; // @[TensorUtil.scala 352:11:@2246.4]
  assign io_stride = _T_176 & _T_181; // @[TensorUtil.scala 347:13:@2232.4]
  assign io_split = _T_173 & _T_184; // @[TensorUtil.scala 348:12:@2233.4]
  assign io_addr = caddr; // @[TensorUtil.scala 350:11:@2236.4]
  assign io_len = len; // @[TensorUtil.scala 351:10:@2237.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  caddr = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  baddr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  len = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  xcnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xrem = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ycnt = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  xfer_bytes = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    caddr <= _GEN_25[31:0];
    baddr <= _GEN_26[31:0];
    len <= _GEN_13[7:0];
    if (io_xinit) begin
      xcnt <= 8'h0;
    end else begin
      if (io_xupdate) begin
        xcnt <= _T_217;
      end
    end
    xrem <= _GEN_14[15:0];
    if (io_start) begin
      ycnt <= 16'h0;
    end else begin
      if (_T_219) begin
        ycnt <= _T_222;
      end
    end
    if (io_start) begin
      xfer_bytes <= {{20'd0}, xfer_init_bytes};
    end else begin
      if (_T_194) begin
        xfer_bytes <= {{20'd0}, xfer_stride_bytes};
      end else begin
        if (_T_204) begin
          xfer_bytes <= {{20'd0}, xfer_split_bytes};
        end
      end
    end
  end
endmodule
module TensorPadCtrl_4( // @[:@2248.2]
  input          clock, // @[:@2249.4]
  input          reset, // @[:@2250.4]
  input          io_start, // @[:@2251.4]
  output         io_done, // @[:@2251.4]
  input  [127:0] io_inst // @[:@2251.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@2276.4]
  wire [3:0] dec_ypad_0; // @[TensorUtil.scala 173:29:@2280.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@2284.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@2286.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@2288.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@2289.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@2290.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@2291.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@2292.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@2292.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@2293.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@2294.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@2294.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@2295.4]
  wire [20:0] _GEN_12; // @[TensorUtil.scala 182:46:@2296.4]
  wire [20:0] _T_39; // @[TensorUtil.scala 182:46:@2296.4]
  wire [21:0] _T_41; // @[TensorUtil.scala 182:71:@2297.4]
  wire [21:0] _T_42; // @[TensorUtil.scala 182:71:@2298.4]
  wire [20:0] xval; // @[TensorUtil.scala 182:71:@2299.4]
  wire  _T_44; // @[TensorUtil.scala 190:22:@2300.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 190:42:@2301.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 190:42:@2302.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 190:42:@2303.4]
  wire [3:0] yval; // @[TensorUtil.scala 190:10:@2304.4]
  reg  state; // @[TensorUtil.scala 197:22:@2305.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@2306.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@2308.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@2315.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@2316.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@2317.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@2318.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@2314.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@2307.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@2322.4]
  wire [20:0] _GEN_4; // @[TensorUtil.scala 212:25:@2323.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@2329.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@2336.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@2337.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@2335.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@2341.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@2342.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@2349.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@2351.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@2352.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@2350.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@2357.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@2276.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorUtil.scala 173:29:@2280.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@2284.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@2286.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@2292.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@2292.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@2293.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@2294.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@2294.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@2295.4]
  assign _GEN_12 = {{5'd0}, _T_38}; // @[TensorUtil.scala 182:46:@2296.4]
  assign _T_39 = _GEN_12 << 5; // @[TensorUtil.scala 182:46:@2296.4]
  assign _T_41 = _T_39 - 21'h1; // @[TensorUtil.scala 182:71:@2297.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@2298.4]
  assign xval = _T_42[20:0]; // @[TensorUtil.scala 182:71:@2299.4]
  assign _T_44 = dec_ypad_0 != 4'h0; // @[TensorUtil.scala 190:22:@2300.4]
  assign _T_46 = dec_ypad_0 - 4'h1; // @[TensorUtil.scala 190:42:@2301.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 190:42:@2302.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 190:42:@2303.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 190:10:@2304.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@2306.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@2308.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@2315.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@2316.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@2317.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@2318.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@2314.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@2307.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@2322.4]
  assign _GEN_4 = _T_56 ? xval : {{5'd0}, xmax}; // @[TensorUtil.scala 212:25:@2323.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@2329.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2336.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2337.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@2335.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@2341.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@2342.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@2349.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@2351.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@2352.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@2350.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@2357.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@2360.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_5( // @[:@2362.2]
  input          clock, // @[:@2363.4]
  input          reset, // @[:@2364.4]
  input          io_start, // @[:@2365.4]
  output         io_done, // @[:@2365.4]
  input  [127:0] io_inst // @[:@2365.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@2390.4]
  wire [3:0] dec_ypad_1; // @[TensorUtil.scala 173:29:@2396.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@2398.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@2400.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@2402.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@2403.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@2404.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@2405.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@2406.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@2406.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@2407.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@2408.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@2408.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@2409.4]
  wire [20:0] _GEN_12; // @[TensorUtil.scala 182:46:@2410.4]
  wire [20:0] _T_39; // @[TensorUtil.scala 182:46:@2410.4]
  wire [21:0] _T_41; // @[TensorUtil.scala 182:71:@2411.4]
  wire [21:0] _T_42; // @[TensorUtil.scala 182:71:@2412.4]
  wire [20:0] xval; // @[TensorUtil.scala 182:71:@2413.4]
  wire  _T_44; // @[TensorUtil.scala 192:22:@2414.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 192:42:@2415.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 192:42:@2416.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 192:42:@2417.4]
  wire [3:0] yval; // @[TensorUtil.scala 192:10:@2418.4]
  reg  state; // @[TensorUtil.scala 197:22:@2419.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@2420.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@2422.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@2429.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@2430.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@2431.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@2432.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@2428.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@2421.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@2436.4]
  wire [20:0] _GEN_4; // @[TensorUtil.scala 212:25:@2437.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@2443.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@2450.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@2451.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@2449.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@2455.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@2456.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@2463.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@2465.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@2466.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@2464.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@2471.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@2390.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorUtil.scala 173:29:@2396.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@2398.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@2400.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@2406.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@2406.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@2407.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@2408.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@2408.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@2409.4]
  assign _GEN_12 = {{5'd0}, _T_38}; // @[TensorUtil.scala 182:46:@2410.4]
  assign _T_39 = _GEN_12 << 5; // @[TensorUtil.scala 182:46:@2410.4]
  assign _T_41 = _T_39 - 21'h1; // @[TensorUtil.scala 182:71:@2411.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@2412.4]
  assign xval = _T_42[20:0]; // @[TensorUtil.scala 182:71:@2413.4]
  assign _T_44 = dec_ypad_1 != 4'h0; // @[TensorUtil.scala 192:22:@2414.4]
  assign _T_46 = dec_ypad_1 - 4'h1; // @[TensorUtil.scala 192:42:@2415.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 192:42:@2416.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 192:42:@2417.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 192:10:@2418.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@2420.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@2422.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@2429.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@2430.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@2431.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@2432.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@2428.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@2421.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@2436.4]
  assign _GEN_4 = _T_56 ? xval : {{5'd0}, xmax}; // @[TensorUtil.scala 212:25:@2437.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@2443.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2450.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2451.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@2449.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@2455.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@2456.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@2463.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@2465.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@2466.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@2464.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@2471.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@2474.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_6( // @[:@2476.2]
  input          clock, // @[:@2477.4]
  input          reset, // @[:@2478.4]
  input          io_start, // @[:@2479.4]
  output         io_done, // @[:@2479.4]
  input  [127:0] io_inst // @[:@2479.4]
);
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@2512.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@2516.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@2518.4]
  reg [31:0] _RAND_1;
  wire [8:0] _GEN_10; // @[TensorUtil.scala 184:19:@2520.4]
  wire [8:0] _T_35; // @[TensorUtil.scala 184:19:@2520.4]
  wire [9:0] _T_37; // @[TensorUtil.scala 184:44:@2521.4]
  wire [9:0] _T_38; // @[TensorUtil.scala 184:44:@2522.4]
  wire [8:0] xval; // @[TensorUtil.scala 184:44:@2523.4]
  reg  state; // @[TensorUtil.scala 197:22:@2524.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@2525.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@2527.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@2535.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@2537.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@2533.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@2526.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@2541.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@2548.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@2555.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@2556.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@2554.6]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@2512.4]
  assign _GEN_10 = {{5'd0}, dec_xpad_0}; // @[TensorUtil.scala 184:19:@2520.4]
  assign _T_35 = _GEN_10 << 5; // @[TensorUtil.scala 184:19:@2520.4]
  assign _T_37 = _T_35 - 9'h1; // @[TensorUtil.scala 184:44:@2521.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 184:44:@2522.4]
  assign xval = _T_38[8:0]; // @[TensorUtil.scala 184:44:@2523.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@2525.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@2527.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@2535.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@2537.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@2533.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@2526.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@2541.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@2548.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2555.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2556.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@2554.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@2579.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{7'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_7( // @[:@2581.2]
  input          clock, // @[:@2582.4]
  input          reset, // @[:@2583.4]
  input          io_start, // @[:@2584.4]
  output         io_done, // @[:@2584.4]
  input  [127:0] io_inst // @[:@2584.4]
);
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@2619.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@2621.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@2623.4]
  reg [31:0] _RAND_1;
  wire [8:0] _GEN_10; // @[TensorUtil.scala 186:19:@2625.4]
  wire [8:0] _T_35; // @[TensorUtil.scala 186:19:@2625.4]
  wire [9:0] _T_37; // @[TensorUtil.scala 186:44:@2626.4]
  wire [9:0] _T_38; // @[TensorUtil.scala 186:44:@2627.4]
  wire [8:0] xval; // @[TensorUtil.scala 186:44:@2628.4]
  reg  state; // @[TensorUtil.scala 197:22:@2629.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@2630.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@2632.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@2640.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@2642.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@2638.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@2631.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@2646.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@2653.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@2660.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@2661.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@2659.6]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@2619.4]
  assign _GEN_10 = {{5'd0}, dec_xpad_1}; // @[TensorUtil.scala 186:19:@2625.4]
  assign _T_35 = _GEN_10 << 5; // @[TensorUtil.scala 186:19:@2625.4]
  assign _T_37 = _T_35 - 9'h1; // @[TensorUtil.scala 186:44:@2626.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 186:44:@2627.4]
  assign xval = _T_38[8:0]; // @[TensorUtil.scala 186:44:@2628.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@2630.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@2632.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@2640.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@2642.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@2638.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@2631.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@2646.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@2653.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2660.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2661.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@2659.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@2684.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{7'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorLoad_1( // @[:@2686.2]
  input          clock, // @[:@2687.4]
  input          reset, // @[:@2688.4]
  input          io_start, // @[:@2689.4]
  output         io_done, // @[:@2689.4]
  input  [127:0] io_inst, // @[:@2689.4]
  input  [31:0]  io_baddr, // @[:@2689.4]
  input          io_vme_rd_cmd_ready, // @[:@2689.4]
  output         io_vme_rd_cmd_valid, // @[:@2689.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@2689.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@2689.4]
  output         io_vme_rd_data_ready, // @[:@2689.4]
  input          io_vme_rd_data_valid, // @[:@2689.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@2689.4]
  input          io_tensor_rd_idx_valid, // @[:@2689.4]
  input  [9:0]   io_tensor_rd_idx_bits, // @[:@2689.4]
  output         io_tensor_rd_data_valid, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_0_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_1_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_2_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_3_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_4_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_5_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_6_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_7_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_8_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_9_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_10_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_11_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_12_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_13_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_14_15, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_0, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_1, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_2, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_3, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_4, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_5, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_6, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_7, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_8, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_9, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_10, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_11, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_12, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_13, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_14, // @[:@2689.4]
  output [7:0]   io_tensor_rd_data_bits_15_15 // @[:@2689.4]
);
  wire  dataCtrl_clock; // @[TensorLoad.scala 52:24:@2726.4]
  wire  dataCtrl_io_start; // @[TensorLoad.scala 52:24:@2726.4]
  wire  dataCtrl_io_done; // @[TensorLoad.scala 52:24:@2726.4]
  wire [127:0] dataCtrl_io_inst; // @[TensorLoad.scala 52:24:@2726.4]
  wire [31:0] dataCtrl_io_baddr; // @[TensorLoad.scala 52:24:@2726.4]
  wire  dataCtrl_io_xinit; // @[TensorLoad.scala 52:24:@2726.4]
  wire  dataCtrl_io_xupdate; // @[TensorLoad.scala 52:24:@2726.4]
  wire  dataCtrl_io_yupdate; // @[TensorLoad.scala 52:24:@2726.4]
  wire  dataCtrl_io_stride; // @[TensorLoad.scala 52:24:@2726.4]
  wire  dataCtrl_io_split; // @[TensorLoad.scala 52:24:@2726.4]
  wire [31:0] dataCtrl_io_addr; // @[TensorLoad.scala 52:24:@2726.4]
  wire [7:0] dataCtrl_io_len; // @[TensorLoad.scala 52:24:@2726.4]
  wire  yPadCtrl0_clock; // @[TensorLoad.scala 55:25:@2730.4]
  wire  yPadCtrl0_reset; // @[TensorLoad.scala 55:25:@2730.4]
  wire  yPadCtrl0_io_start; // @[TensorLoad.scala 55:25:@2730.4]
  wire  yPadCtrl0_io_done; // @[TensorLoad.scala 55:25:@2730.4]
  wire [127:0] yPadCtrl0_io_inst; // @[TensorLoad.scala 55:25:@2730.4]
  wire  yPadCtrl1_clock; // @[TensorLoad.scala 56:25:@2733.4]
  wire  yPadCtrl1_reset; // @[TensorLoad.scala 56:25:@2733.4]
  wire  yPadCtrl1_io_start; // @[TensorLoad.scala 56:25:@2733.4]
  wire  yPadCtrl1_io_done; // @[TensorLoad.scala 56:25:@2733.4]
  wire [127:0] yPadCtrl1_io_inst; // @[TensorLoad.scala 56:25:@2733.4]
  wire  xPadCtrl0_clock; // @[TensorLoad.scala 57:25:@2736.4]
  wire  xPadCtrl0_reset; // @[TensorLoad.scala 57:25:@2736.4]
  wire  xPadCtrl0_io_start; // @[TensorLoad.scala 57:25:@2736.4]
  wire  xPadCtrl0_io_done; // @[TensorLoad.scala 57:25:@2736.4]
  wire [127:0] xPadCtrl0_io_inst; // @[TensorLoad.scala 57:25:@2736.4]
  wire  xPadCtrl1_clock; // @[TensorLoad.scala 58:25:@2739.4]
  wire  xPadCtrl1_reset; // @[TensorLoad.scala 58:25:@2739.4]
  wire  xPadCtrl1_io_start; // @[TensorLoad.scala 58:25:@2739.4]
  wire  xPadCtrl1_io_done; // @[TensorLoad.scala 58:25:@2739.4]
  wire [127:0] xPadCtrl1_io_inst; // @[TensorLoad.scala 58:25:@2739.4]
  reg [63:0] tensorFile_0_0 [0:1023]; // @[TensorLoad.scala 222:16:@3009.4]
  reg [63:0] _RAND_0;
  wire [63:0] tensorFile_0_0_rdata_0_data; // @[TensorLoad.scala 222:16:@3009.4]
  wire [9:0] tensorFile_0_0_rdata_0_addr; // @[TensorLoad.scala 222:16:@3009.4]
  wire [63:0] tensorFile_0_0__T_4976_data; // @[TensorLoad.scala 222:16:@3009.4]
  wire [9:0] tensorFile_0_0__T_4976_addr; // @[TensorLoad.scala 222:16:@3009.4]
  wire  tensorFile_0_0__T_4976_mask; // @[TensorLoad.scala 222:16:@3009.4]
  wire  tensorFile_0_0__T_4976_en; // @[TensorLoad.scala 222:16:@3009.4]
  reg [63:0] tensorFile_0_1 [0:1023]; // @[TensorLoad.scala 222:16:@3009.4]
  reg [63:0] _RAND_1;
  wire [63:0] tensorFile_0_1_rdata_0_data; // @[TensorLoad.scala 222:16:@3009.4]
  wire [9:0] tensorFile_0_1_rdata_0_addr; // @[TensorLoad.scala 222:16:@3009.4]
  wire [63:0] tensorFile_0_1__T_4976_data; // @[TensorLoad.scala 222:16:@3009.4]
  wire [9:0] tensorFile_0_1__T_4976_addr; // @[TensorLoad.scala 222:16:@3009.4]
  wire  tensorFile_0_1__T_4976_mask; // @[TensorLoad.scala 222:16:@3009.4]
  wire  tensorFile_0_1__T_4976_en; // @[TensorLoad.scala 222:16:@3009.4]
  reg [63:0] tensorFile_1_0 [0:1023]; // @[TensorLoad.scala 222:16:@3010.4]
  reg [63:0] _RAND_2;
  wire [63:0] tensorFile_1_0_rdata_1_data; // @[TensorLoad.scala 222:16:@3010.4]
  wire [9:0] tensorFile_1_0_rdata_1_addr; // @[TensorLoad.scala 222:16:@3010.4]
  wire [63:0] tensorFile_1_0__T_5063_data; // @[TensorLoad.scala 222:16:@3010.4]
  wire [9:0] tensorFile_1_0__T_5063_addr; // @[TensorLoad.scala 222:16:@3010.4]
  wire  tensorFile_1_0__T_5063_mask; // @[TensorLoad.scala 222:16:@3010.4]
  wire  tensorFile_1_0__T_5063_en; // @[TensorLoad.scala 222:16:@3010.4]
  reg [63:0] tensorFile_1_1 [0:1023]; // @[TensorLoad.scala 222:16:@3010.4]
  reg [63:0] _RAND_3;
  wire [63:0] tensorFile_1_1_rdata_1_data; // @[TensorLoad.scala 222:16:@3010.4]
  wire [9:0] tensorFile_1_1_rdata_1_addr; // @[TensorLoad.scala 222:16:@3010.4]
  wire [63:0] tensorFile_1_1__T_5063_data; // @[TensorLoad.scala 222:16:@3010.4]
  wire [9:0] tensorFile_1_1__T_5063_addr; // @[TensorLoad.scala 222:16:@3010.4]
  wire  tensorFile_1_1__T_5063_mask; // @[TensorLoad.scala 222:16:@3010.4]
  wire  tensorFile_1_1__T_5063_en; // @[TensorLoad.scala 222:16:@3010.4]
  reg [63:0] tensorFile_2_0 [0:1023]; // @[TensorLoad.scala 222:16:@3011.4]
  reg [63:0] _RAND_4;
  wire [63:0] tensorFile_2_0_rdata_2_data; // @[TensorLoad.scala 222:16:@3011.4]
  wire [9:0] tensorFile_2_0_rdata_2_addr; // @[TensorLoad.scala 222:16:@3011.4]
  wire [63:0] tensorFile_2_0__T_5150_data; // @[TensorLoad.scala 222:16:@3011.4]
  wire [9:0] tensorFile_2_0__T_5150_addr; // @[TensorLoad.scala 222:16:@3011.4]
  wire  tensorFile_2_0__T_5150_mask; // @[TensorLoad.scala 222:16:@3011.4]
  wire  tensorFile_2_0__T_5150_en; // @[TensorLoad.scala 222:16:@3011.4]
  reg [63:0] tensorFile_2_1 [0:1023]; // @[TensorLoad.scala 222:16:@3011.4]
  reg [63:0] _RAND_5;
  wire [63:0] tensorFile_2_1_rdata_2_data; // @[TensorLoad.scala 222:16:@3011.4]
  wire [9:0] tensorFile_2_1_rdata_2_addr; // @[TensorLoad.scala 222:16:@3011.4]
  wire [63:0] tensorFile_2_1__T_5150_data; // @[TensorLoad.scala 222:16:@3011.4]
  wire [9:0] tensorFile_2_1__T_5150_addr; // @[TensorLoad.scala 222:16:@3011.4]
  wire  tensorFile_2_1__T_5150_mask; // @[TensorLoad.scala 222:16:@3011.4]
  wire  tensorFile_2_1__T_5150_en; // @[TensorLoad.scala 222:16:@3011.4]
  reg [63:0] tensorFile_3_0 [0:1023]; // @[TensorLoad.scala 222:16:@3012.4]
  reg [63:0] _RAND_6;
  wire [63:0] tensorFile_3_0_rdata_3_data; // @[TensorLoad.scala 222:16:@3012.4]
  wire [9:0] tensorFile_3_0_rdata_3_addr; // @[TensorLoad.scala 222:16:@3012.4]
  wire [63:0] tensorFile_3_0__T_5237_data; // @[TensorLoad.scala 222:16:@3012.4]
  wire [9:0] tensorFile_3_0__T_5237_addr; // @[TensorLoad.scala 222:16:@3012.4]
  wire  tensorFile_3_0__T_5237_mask; // @[TensorLoad.scala 222:16:@3012.4]
  wire  tensorFile_3_0__T_5237_en; // @[TensorLoad.scala 222:16:@3012.4]
  reg [63:0] tensorFile_3_1 [0:1023]; // @[TensorLoad.scala 222:16:@3012.4]
  reg [63:0] _RAND_7;
  wire [63:0] tensorFile_3_1_rdata_3_data; // @[TensorLoad.scala 222:16:@3012.4]
  wire [9:0] tensorFile_3_1_rdata_3_addr; // @[TensorLoad.scala 222:16:@3012.4]
  wire [63:0] tensorFile_3_1__T_5237_data; // @[TensorLoad.scala 222:16:@3012.4]
  wire [9:0] tensorFile_3_1__T_5237_addr; // @[TensorLoad.scala 222:16:@3012.4]
  wire  tensorFile_3_1__T_5237_mask; // @[TensorLoad.scala 222:16:@3012.4]
  wire  tensorFile_3_1__T_5237_en; // @[TensorLoad.scala 222:16:@3012.4]
  reg [63:0] tensorFile_4_0 [0:1023]; // @[TensorLoad.scala 222:16:@3013.4]
  reg [63:0] _RAND_8;
  wire [63:0] tensorFile_4_0_rdata_4_data; // @[TensorLoad.scala 222:16:@3013.4]
  wire [9:0] tensorFile_4_0_rdata_4_addr; // @[TensorLoad.scala 222:16:@3013.4]
  wire [63:0] tensorFile_4_0__T_5324_data; // @[TensorLoad.scala 222:16:@3013.4]
  wire [9:0] tensorFile_4_0__T_5324_addr; // @[TensorLoad.scala 222:16:@3013.4]
  wire  tensorFile_4_0__T_5324_mask; // @[TensorLoad.scala 222:16:@3013.4]
  wire  tensorFile_4_0__T_5324_en; // @[TensorLoad.scala 222:16:@3013.4]
  reg [63:0] tensorFile_4_1 [0:1023]; // @[TensorLoad.scala 222:16:@3013.4]
  reg [63:0] _RAND_9;
  wire [63:0] tensorFile_4_1_rdata_4_data; // @[TensorLoad.scala 222:16:@3013.4]
  wire [9:0] tensorFile_4_1_rdata_4_addr; // @[TensorLoad.scala 222:16:@3013.4]
  wire [63:0] tensorFile_4_1__T_5324_data; // @[TensorLoad.scala 222:16:@3013.4]
  wire [9:0] tensorFile_4_1__T_5324_addr; // @[TensorLoad.scala 222:16:@3013.4]
  wire  tensorFile_4_1__T_5324_mask; // @[TensorLoad.scala 222:16:@3013.4]
  wire  tensorFile_4_1__T_5324_en; // @[TensorLoad.scala 222:16:@3013.4]
  reg [63:0] tensorFile_5_0 [0:1023]; // @[TensorLoad.scala 222:16:@3014.4]
  reg [63:0] _RAND_10;
  wire [63:0] tensorFile_5_0_rdata_5_data; // @[TensorLoad.scala 222:16:@3014.4]
  wire [9:0] tensorFile_5_0_rdata_5_addr; // @[TensorLoad.scala 222:16:@3014.4]
  wire [63:0] tensorFile_5_0__T_5411_data; // @[TensorLoad.scala 222:16:@3014.4]
  wire [9:0] tensorFile_5_0__T_5411_addr; // @[TensorLoad.scala 222:16:@3014.4]
  wire  tensorFile_5_0__T_5411_mask; // @[TensorLoad.scala 222:16:@3014.4]
  wire  tensorFile_5_0__T_5411_en; // @[TensorLoad.scala 222:16:@3014.4]
  reg [63:0] tensorFile_5_1 [0:1023]; // @[TensorLoad.scala 222:16:@3014.4]
  reg [63:0] _RAND_11;
  wire [63:0] tensorFile_5_1_rdata_5_data; // @[TensorLoad.scala 222:16:@3014.4]
  wire [9:0] tensorFile_5_1_rdata_5_addr; // @[TensorLoad.scala 222:16:@3014.4]
  wire [63:0] tensorFile_5_1__T_5411_data; // @[TensorLoad.scala 222:16:@3014.4]
  wire [9:0] tensorFile_5_1__T_5411_addr; // @[TensorLoad.scala 222:16:@3014.4]
  wire  tensorFile_5_1__T_5411_mask; // @[TensorLoad.scala 222:16:@3014.4]
  wire  tensorFile_5_1__T_5411_en; // @[TensorLoad.scala 222:16:@3014.4]
  reg [63:0] tensorFile_6_0 [0:1023]; // @[TensorLoad.scala 222:16:@3015.4]
  reg [63:0] _RAND_12;
  wire [63:0] tensorFile_6_0_rdata_6_data; // @[TensorLoad.scala 222:16:@3015.4]
  wire [9:0] tensorFile_6_0_rdata_6_addr; // @[TensorLoad.scala 222:16:@3015.4]
  wire [63:0] tensorFile_6_0__T_5498_data; // @[TensorLoad.scala 222:16:@3015.4]
  wire [9:0] tensorFile_6_0__T_5498_addr; // @[TensorLoad.scala 222:16:@3015.4]
  wire  tensorFile_6_0__T_5498_mask; // @[TensorLoad.scala 222:16:@3015.4]
  wire  tensorFile_6_0__T_5498_en; // @[TensorLoad.scala 222:16:@3015.4]
  reg [63:0] tensorFile_6_1 [0:1023]; // @[TensorLoad.scala 222:16:@3015.4]
  reg [63:0] _RAND_13;
  wire [63:0] tensorFile_6_1_rdata_6_data; // @[TensorLoad.scala 222:16:@3015.4]
  wire [9:0] tensorFile_6_1_rdata_6_addr; // @[TensorLoad.scala 222:16:@3015.4]
  wire [63:0] tensorFile_6_1__T_5498_data; // @[TensorLoad.scala 222:16:@3015.4]
  wire [9:0] tensorFile_6_1__T_5498_addr; // @[TensorLoad.scala 222:16:@3015.4]
  wire  tensorFile_6_1__T_5498_mask; // @[TensorLoad.scala 222:16:@3015.4]
  wire  tensorFile_6_1__T_5498_en; // @[TensorLoad.scala 222:16:@3015.4]
  reg [63:0] tensorFile_7_0 [0:1023]; // @[TensorLoad.scala 222:16:@3016.4]
  reg [63:0] _RAND_14;
  wire [63:0] tensorFile_7_0_rdata_7_data; // @[TensorLoad.scala 222:16:@3016.4]
  wire [9:0] tensorFile_7_0_rdata_7_addr; // @[TensorLoad.scala 222:16:@3016.4]
  wire [63:0] tensorFile_7_0__T_5585_data; // @[TensorLoad.scala 222:16:@3016.4]
  wire [9:0] tensorFile_7_0__T_5585_addr; // @[TensorLoad.scala 222:16:@3016.4]
  wire  tensorFile_7_0__T_5585_mask; // @[TensorLoad.scala 222:16:@3016.4]
  wire  tensorFile_7_0__T_5585_en; // @[TensorLoad.scala 222:16:@3016.4]
  reg [63:0] tensorFile_7_1 [0:1023]; // @[TensorLoad.scala 222:16:@3016.4]
  reg [63:0] _RAND_15;
  wire [63:0] tensorFile_7_1_rdata_7_data; // @[TensorLoad.scala 222:16:@3016.4]
  wire [9:0] tensorFile_7_1_rdata_7_addr; // @[TensorLoad.scala 222:16:@3016.4]
  wire [63:0] tensorFile_7_1__T_5585_data; // @[TensorLoad.scala 222:16:@3016.4]
  wire [9:0] tensorFile_7_1__T_5585_addr; // @[TensorLoad.scala 222:16:@3016.4]
  wire  tensorFile_7_1__T_5585_mask; // @[TensorLoad.scala 222:16:@3016.4]
  wire  tensorFile_7_1__T_5585_en; // @[TensorLoad.scala 222:16:@3016.4]
  reg [63:0] tensorFile_8_0 [0:1023]; // @[TensorLoad.scala 222:16:@3017.4]
  reg [63:0] _RAND_16;
  wire [63:0] tensorFile_8_0_rdata_8_data; // @[TensorLoad.scala 222:16:@3017.4]
  wire [9:0] tensorFile_8_0_rdata_8_addr; // @[TensorLoad.scala 222:16:@3017.4]
  wire [63:0] tensorFile_8_0__T_5672_data; // @[TensorLoad.scala 222:16:@3017.4]
  wire [9:0] tensorFile_8_0__T_5672_addr; // @[TensorLoad.scala 222:16:@3017.4]
  wire  tensorFile_8_0__T_5672_mask; // @[TensorLoad.scala 222:16:@3017.4]
  wire  tensorFile_8_0__T_5672_en; // @[TensorLoad.scala 222:16:@3017.4]
  reg [63:0] tensorFile_8_1 [0:1023]; // @[TensorLoad.scala 222:16:@3017.4]
  reg [63:0] _RAND_17;
  wire [63:0] tensorFile_8_1_rdata_8_data; // @[TensorLoad.scala 222:16:@3017.4]
  wire [9:0] tensorFile_8_1_rdata_8_addr; // @[TensorLoad.scala 222:16:@3017.4]
  wire [63:0] tensorFile_8_1__T_5672_data; // @[TensorLoad.scala 222:16:@3017.4]
  wire [9:0] tensorFile_8_1__T_5672_addr; // @[TensorLoad.scala 222:16:@3017.4]
  wire  tensorFile_8_1__T_5672_mask; // @[TensorLoad.scala 222:16:@3017.4]
  wire  tensorFile_8_1__T_5672_en; // @[TensorLoad.scala 222:16:@3017.4]
  reg [63:0] tensorFile_9_0 [0:1023]; // @[TensorLoad.scala 222:16:@3018.4]
  reg [63:0] _RAND_18;
  wire [63:0] tensorFile_9_0_rdata_9_data; // @[TensorLoad.scala 222:16:@3018.4]
  wire [9:0] tensorFile_9_0_rdata_9_addr; // @[TensorLoad.scala 222:16:@3018.4]
  wire [63:0] tensorFile_9_0__T_5759_data; // @[TensorLoad.scala 222:16:@3018.4]
  wire [9:0] tensorFile_9_0__T_5759_addr; // @[TensorLoad.scala 222:16:@3018.4]
  wire  tensorFile_9_0__T_5759_mask; // @[TensorLoad.scala 222:16:@3018.4]
  wire  tensorFile_9_0__T_5759_en; // @[TensorLoad.scala 222:16:@3018.4]
  reg [63:0] tensorFile_9_1 [0:1023]; // @[TensorLoad.scala 222:16:@3018.4]
  reg [63:0] _RAND_19;
  wire [63:0] tensorFile_9_1_rdata_9_data; // @[TensorLoad.scala 222:16:@3018.4]
  wire [9:0] tensorFile_9_1_rdata_9_addr; // @[TensorLoad.scala 222:16:@3018.4]
  wire [63:0] tensorFile_9_1__T_5759_data; // @[TensorLoad.scala 222:16:@3018.4]
  wire [9:0] tensorFile_9_1__T_5759_addr; // @[TensorLoad.scala 222:16:@3018.4]
  wire  tensorFile_9_1__T_5759_mask; // @[TensorLoad.scala 222:16:@3018.4]
  wire  tensorFile_9_1__T_5759_en; // @[TensorLoad.scala 222:16:@3018.4]
  reg [63:0] tensorFile_10_0 [0:1023]; // @[TensorLoad.scala 222:16:@3019.4]
  reg [63:0] _RAND_20;
  wire [63:0] tensorFile_10_0_rdata_10_data; // @[TensorLoad.scala 222:16:@3019.4]
  wire [9:0] tensorFile_10_0_rdata_10_addr; // @[TensorLoad.scala 222:16:@3019.4]
  wire [63:0] tensorFile_10_0__T_5846_data; // @[TensorLoad.scala 222:16:@3019.4]
  wire [9:0] tensorFile_10_0__T_5846_addr; // @[TensorLoad.scala 222:16:@3019.4]
  wire  tensorFile_10_0__T_5846_mask; // @[TensorLoad.scala 222:16:@3019.4]
  wire  tensorFile_10_0__T_5846_en; // @[TensorLoad.scala 222:16:@3019.4]
  reg [63:0] tensorFile_10_1 [0:1023]; // @[TensorLoad.scala 222:16:@3019.4]
  reg [63:0] _RAND_21;
  wire [63:0] tensorFile_10_1_rdata_10_data; // @[TensorLoad.scala 222:16:@3019.4]
  wire [9:0] tensorFile_10_1_rdata_10_addr; // @[TensorLoad.scala 222:16:@3019.4]
  wire [63:0] tensorFile_10_1__T_5846_data; // @[TensorLoad.scala 222:16:@3019.4]
  wire [9:0] tensorFile_10_1__T_5846_addr; // @[TensorLoad.scala 222:16:@3019.4]
  wire  tensorFile_10_1__T_5846_mask; // @[TensorLoad.scala 222:16:@3019.4]
  wire  tensorFile_10_1__T_5846_en; // @[TensorLoad.scala 222:16:@3019.4]
  reg [63:0] tensorFile_11_0 [0:1023]; // @[TensorLoad.scala 222:16:@3020.4]
  reg [63:0] _RAND_22;
  wire [63:0] tensorFile_11_0_rdata_11_data; // @[TensorLoad.scala 222:16:@3020.4]
  wire [9:0] tensorFile_11_0_rdata_11_addr; // @[TensorLoad.scala 222:16:@3020.4]
  wire [63:0] tensorFile_11_0__T_5933_data; // @[TensorLoad.scala 222:16:@3020.4]
  wire [9:0] tensorFile_11_0__T_5933_addr; // @[TensorLoad.scala 222:16:@3020.4]
  wire  tensorFile_11_0__T_5933_mask; // @[TensorLoad.scala 222:16:@3020.4]
  wire  tensorFile_11_0__T_5933_en; // @[TensorLoad.scala 222:16:@3020.4]
  reg [63:0] tensorFile_11_1 [0:1023]; // @[TensorLoad.scala 222:16:@3020.4]
  reg [63:0] _RAND_23;
  wire [63:0] tensorFile_11_1_rdata_11_data; // @[TensorLoad.scala 222:16:@3020.4]
  wire [9:0] tensorFile_11_1_rdata_11_addr; // @[TensorLoad.scala 222:16:@3020.4]
  wire [63:0] tensorFile_11_1__T_5933_data; // @[TensorLoad.scala 222:16:@3020.4]
  wire [9:0] tensorFile_11_1__T_5933_addr; // @[TensorLoad.scala 222:16:@3020.4]
  wire  tensorFile_11_1__T_5933_mask; // @[TensorLoad.scala 222:16:@3020.4]
  wire  tensorFile_11_1__T_5933_en; // @[TensorLoad.scala 222:16:@3020.4]
  reg [63:0] tensorFile_12_0 [0:1023]; // @[TensorLoad.scala 222:16:@3021.4]
  reg [63:0] _RAND_24;
  wire [63:0] tensorFile_12_0_rdata_12_data; // @[TensorLoad.scala 222:16:@3021.4]
  wire [9:0] tensorFile_12_0_rdata_12_addr; // @[TensorLoad.scala 222:16:@3021.4]
  wire [63:0] tensorFile_12_0__T_6020_data; // @[TensorLoad.scala 222:16:@3021.4]
  wire [9:0] tensorFile_12_0__T_6020_addr; // @[TensorLoad.scala 222:16:@3021.4]
  wire  tensorFile_12_0__T_6020_mask; // @[TensorLoad.scala 222:16:@3021.4]
  wire  tensorFile_12_0__T_6020_en; // @[TensorLoad.scala 222:16:@3021.4]
  reg [63:0] tensorFile_12_1 [0:1023]; // @[TensorLoad.scala 222:16:@3021.4]
  reg [63:0] _RAND_25;
  wire [63:0] tensorFile_12_1_rdata_12_data; // @[TensorLoad.scala 222:16:@3021.4]
  wire [9:0] tensorFile_12_1_rdata_12_addr; // @[TensorLoad.scala 222:16:@3021.4]
  wire [63:0] tensorFile_12_1__T_6020_data; // @[TensorLoad.scala 222:16:@3021.4]
  wire [9:0] tensorFile_12_1__T_6020_addr; // @[TensorLoad.scala 222:16:@3021.4]
  wire  tensorFile_12_1__T_6020_mask; // @[TensorLoad.scala 222:16:@3021.4]
  wire  tensorFile_12_1__T_6020_en; // @[TensorLoad.scala 222:16:@3021.4]
  reg [63:0] tensorFile_13_0 [0:1023]; // @[TensorLoad.scala 222:16:@3022.4]
  reg [63:0] _RAND_26;
  wire [63:0] tensorFile_13_0_rdata_13_data; // @[TensorLoad.scala 222:16:@3022.4]
  wire [9:0] tensorFile_13_0_rdata_13_addr; // @[TensorLoad.scala 222:16:@3022.4]
  wire [63:0] tensorFile_13_0__T_6107_data; // @[TensorLoad.scala 222:16:@3022.4]
  wire [9:0] tensorFile_13_0__T_6107_addr; // @[TensorLoad.scala 222:16:@3022.4]
  wire  tensorFile_13_0__T_6107_mask; // @[TensorLoad.scala 222:16:@3022.4]
  wire  tensorFile_13_0__T_6107_en; // @[TensorLoad.scala 222:16:@3022.4]
  reg [63:0] tensorFile_13_1 [0:1023]; // @[TensorLoad.scala 222:16:@3022.4]
  reg [63:0] _RAND_27;
  wire [63:0] tensorFile_13_1_rdata_13_data; // @[TensorLoad.scala 222:16:@3022.4]
  wire [9:0] tensorFile_13_1_rdata_13_addr; // @[TensorLoad.scala 222:16:@3022.4]
  wire [63:0] tensorFile_13_1__T_6107_data; // @[TensorLoad.scala 222:16:@3022.4]
  wire [9:0] tensorFile_13_1__T_6107_addr; // @[TensorLoad.scala 222:16:@3022.4]
  wire  tensorFile_13_1__T_6107_mask; // @[TensorLoad.scala 222:16:@3022.4]
  wire  tensorFile_13_1__T_6107_en; // @[TensorLoad.scala 222:16:@3022.4]
  reg [63:0] tensorFile_14_0 [0:1023]; // @[TensorLoad.scala 222:16:@3023.4]
  reg [63:0] _RAND_28;
  wire [63:0] tensorFile_14_0_rdata_14_data; // @[TensorLoad.scala 222:16:@3023.4]
  wire [9:0] tensorFile_14_0_rdata_14_addr; // @[TensorLoad.scala 222:16:@3023.4]
  wire [63:0] tensorFile_14_0__T_6194_data; // @[TensorLoad.scala 222:16:@3023.4]
  wire [9:0] tensorFile_14_0__T_6194_addr; // @[TensorLoad.scala 222:16:@3023.4]
  wire  tensorFile_14_0__T_6194_mask; // @[TensorLoad.scala 222:16:@3023.4]
  wire  tensorFile_14_0__T_6194_en; // @[TensorLoad.scala 222:16:@3023.4]
  reg [63:0] tensorFile_14_1 [0:1023]; // @[TensorLoad.scala 222:16:@3023.4]
  reg [63:0] _RAND_29;
  wire [63:0] tensorFile_14_1_rdata_14_data; // @[TensorLoad.scala 222:16:@3023.4]
  wire [9:0] tensorFile_14_1_rdata_14_addr; // @[TensorLoad.scala 222:16:@3023.4]
  wire [63:0] tensorFile_14_1__T_6194_data; // @[TensorLoad.scala 222:16:@3023.4]
  wire [9:0] tensorFile_14_1__T_6194_addr; // @[TensorLoad.scala 222:16:@3023.4]
  wire  tensorFile_14_1__T_6194_mask; // @[TensorLoad.scala 222:16:@3023.4]
  wire  tensorFile_14_1__T_6194_en; // @[TensorLoad.scala 222:16:@3023.4]
  reg [63:0] tensorFile_15_0 [0:1023]; // @[TensorLoad.scala 222:16:@3024.4]
  reg [63:0] _RAND_30;
  wire [63:0] tensorFile_15_0_rdata_15_data; // @[TensorLoad.scala 222:16:@3024.4]
  wire [9:0] tensorFile_15_0_rdata_15_addr; // @[TensorLoad.scala 222:16:@3024.4]
  wire [63:0] tensorFile_15_0__T_6281_data; // @[TensorLoad.scala 222:16:@3024.4]
  wire [9:0] tensorFile_15_0__T_6281_addr; // @[TensorLoad.scala 222:16:@3024.4]
  wire  tensorFile_15_0__T_6281_mask; // @[TensorLoad.scala 222:16:@3024.4]
  wire  tensorFile_15_0__T_6281_en; // @[TensorLoad.scala 222:16:@3024.4]
  reg [63:0] tensorFile_15_1 [0:1023]; // @[TensorLoad.scala 222:16:@3024.4]
  reg [63:0] _RAND_31;
  wire [63:0] tensorFile_15_1_rdata_15_data; // @[TensorLoad.scala 222:16:@3024.4]
  wire [9:0] tensorFile_15_1_rdata_15_addr; // @[TensorLoad.scala 222:16:@3024.4]
  wire [63:0] tensorFile_15_1__T_6281_data; // @[TensorLoad.scala 222:16:@3024.4]
  wire [9:0] tensorFile_15_1__T_6281_addr; // @[TensorLoad.scala 222:16:@3024.4]
  wire  tensorFile_15_1__T_6281_mask; // @[TensorLoad.scala 222:16:@3024.4]
  wire  tensorFile_15_1__T_6281_en; // @[TensorLoad.scala 222:16:@3024.4]
  wire [15:0] dec_sram_offset; // @[TensorLoad.scala 51:29:@2706.4]
  wire [15:0] dec_xsize; // @[TensorLoad.scala 51:29:@2714.4]
  wire [3:0] dec_ypad_0; // @[TensorLoad.scala 51:29:@2718.4]
  wire [3:0] dec_ypad_1; // @[TensorLoad.scala 51:29:@2720.4]
  wire [3:0] dec_xpad_0; // @[TensorLoad.scala 51:29:@2722.4]
  wire [3:0] dec_xpad_1; // @[TensorLoad.scala 51:29:@2724.4]
  reg  dataCtrlDone; // @[TensorLoad.scala 54:29:@2729.4]
  reg [31:0] _RAND_32;
  reg  tag; // @[TensorLoad.scala 60:16:@2742.4]
  reg [31:0] _RAND_33;
  reg [3:0] set; // @[TensorLoad.scala 61:16:@2743.4]
  reg [31:0] _RAND_34;
  reg [2:0] state; // @[TensorLoad.scala 65:22:@2744.4]
  reg [31:0] _RAND_35;
  wire  _T_4394; // @[Conditional.scala 37:30:@2745.4]
  wire  _T_4396; // @[TensorLoad.scala 71:25:@2748.8]
  wire  _T_4398; // @[TensorLoad.scala 73:31:@2753.10]
  wire [2:0] _GEN_0; // @[TensorLoad.scala 73:40:@2754.10]
  wire [2:0] _GEN_1; // @[TensorLoad.scala 71:34:@2749.8]
  wire [2:0] _GEN_2; // @[TensorLoad.scala 70:22:@2747.6]
  wire  _T_4399; // @[Conditional.scala 37:30:@2763.6]
  wire [2:0] _GEN_4; // @[TensorLoad.scala 81:31:@2765.8]
  wire  _T_4402; // @[Conditional.scala 37:30:@2776.8]
  wire [2:0] _GEN_5; // @[TensorLoad.scala 90:31:@2778.10]
  wire  _T_4403; // @[Conditional.scala 37:30:@2783.10]
  wire [2:0] _GEN_6; // @[TensorLoad.scala 95:33:@2785.12]
  wire  _T_4404; // @[Conditional.scala 37:30:@2790.12]
  wire  _T_4406; // @[TensorLoad.scala 102:27:@2794.18]
  wire  _T_4408; // @[TensorLoad.scala 104:33:@2799.20]
  wire [2:0] _GEN_7; // @[TensorLoad.scala 104:42:@2800.20]
  wire [2:0] _GEN_8; // @[TensorLoad.scala 102:36:@2795.18]
  wire [2:0] _GEN_10; // @[TensorLoad.scala 110:36:@2810.20]
  wire [2:0] _GEN_11; // @[TensorLoad.scala 117:39:@2823.20]
  wire [2:0] _GEN_12; // @[TensorLoad.scala 109:40:@2808.18]
  wire [2:0] _GEN_13; // @[TensorLoad.scala 101:32:@2793.16]
  wire [2:0] _GEN_14; // @[TensorLoad.scala 100:34:@2792.14]
  wire  _T_4413; // @[Conditional.scala 37:30:@2829.14]
  wire [2:0] _GEN_17; // @[TensorLoad.scala 124:28:@2832.18]
  wire [2:0] _GEN_18; // @[TensorLoad.scala 123:31:@2831.16]
  wire  _T_4418; // @[Conditional.scala 37:30:@2853.16]
  wire  _T_4419; // @[TensorLoad.scala 140:30:@2855.18]
  wire [2:0] _GEN_19; // @[TensorLoad.scala 140:47:@2856.18]
  wire [2:0] _GEN_20; // @[Conditional.scala 39:67:@2854.16]
  wire [2:0] _GEN_21; // @[Conditional.scala 39:67:@2830.14]
  wire [2:0] _GEN_22; // @[Conditional.scala 39:67:@2791.12]
  wire [2:0] _GEN_23; // @[Conditional.scala 39:67:@2784.10]
  wire [2:0] _GEN_24; // @[Conditional.scala 39:67:@2777.8]
  wire [2:0] _GEN_25; // @[Conditional.scala 39:67:@2764.6]
  wire [2:0] _GEN_26; // @[Conditional.scala 40:58:@2746.4]
  wire  _T_4420; // @[TensorLoad.scala 147:30:@2860.4]
  wire  _T_4421; // @[TensorLoad.scala 147:40:@2861.4]
  wire  _T_4423; // @[Decoupled.scala 37:37:@2867.4]
  wire  _T_4428; // @[TensorLoad.scala 156:36:@2877.6]
  wire  _GEN_27; // @[TensorLoad.scala 156:57:@2878.6]
  wire  _GEN_28; // @[TensorLoad.scala 154:25:@2872.4]
  wire  _T_4433; // @[TensorLoad.scala 161:44:@2883.4]
  wire  _T_4440; // @[TensorLoad.scala 164:61:@2889.4]
  wire  _T_4441; // @[TensorLoad.scala 164:48:@2890.4]
  wire  _T_4442; // @[TensorLoad.scala 165:14:@2891.4]
  wire  _T_4443; // @[TensorLoad.scala 165:25:@2892.4]
  wire  _T_4444; // @[TensorLoad.scala 165:45:@2893.4]
  wire  _T_4445; // @[TensorLoad.scala 164:70:@2894.4]
  wire  _T_4451; // @[TensorLoad.scala 169:14:@2900.4]
  wire  _T_4452; // @[TensorLoad.scala 169:25:@2901.4]
  wire  _T_4453; // @[TensorLoad.scala 168:35:@2902.4]
  wire  _T_4455; // @[TensorLoad.scala 170:32:@2904.4]
  wire  _T_4456; // @[TensorLoad.scala 170:30:@2905.4]
  wire  _T_4457; // @[TensorLoad.scala 170:46:@2906.4]
  wire  _T_4460; // @[TensorLoad.scala 170:67:@2908.4]
  wire  _T_4461; // @[TensorLoad.scala 169:46:@2909.4]
  wire  _T_4465; // @[TensorLoad.scala 171:45:@2913.4]
  wire  _T_4466; // @[TensorLoad.scala 170:89:@2914.4]
  wire  _T_4471; // @[TensorLoad.scala 173:44:@2919.4]
  wire  _T_4472; // @[TensorLoad.scala 174:28:@2920.4]
  wire  _T_4473; // @[TensorLoad.scala 174:46:@2921.4]
  wire  _T_4476; // @[TensorLoad.scala 174:67:@2923.4]
  wire  _T_4477; // @[TensorLoad.scala 174:25:@2924.4]
  wire  _T_4479; // @[TensorLoad.scala 182:32:@2931.4]
  wire  _T_4482; // @[TensorLoad.scala 190:11:@2938.4]
  wire  _T_4483; // @[TensorLoad.scala 189:36:@2939.4]
  wire  _T_4485; // @[TensorLoad.scala 190:22:@2941.4]
  wire  _T_4486; // @[TensorLoad.scala 192:11:@2942.4]
  wire  isZeroPad; // @[TensorLoad.scala 191:22:@2943.4]
  wire  _T_4489; // @[TensorLoad.scala 194:24:@2946.4]
  wire  _T_4492; // @[TensorLoad.scala 194:46:@2948.4]
  wire  _T_4495; // @[TensorLoad.scala 196:36:@2954.6]
  wire [1:0] _T_4497; // @[TensorLoad.scala 197:16:@2956.8]
  wire  _T_4498; // @[TensorLoad.scala 197:16:@2957.8]
  wire  _GEN_29; // @[TensorLoad.scala 196:50:@2955.6]
  wire  _T_4500; // @[TensorLoad.scala 200:24:@2961.4]
  wire  _T_4502; // @[TensorLoad.scala 200:48:@2962.4]
  wire  _T_4505; // @[TensorLoad.scala 200:76:@2964.4]
  wire  _T_4506; // @[TensorLoad.scala 200:40:@2965.4]
  wire  _T_4512; // @[TensorLoad.scala 202:51:@2973.6]
  wire [4:0] _T_4514; // @[TensorLoad.scala 203:16:@2975.8]
  wire [3:0] _T_4515; // @[TensorLoad.scala 203:16:@2976.8]
  wire [3:0] _GEN_31; // @[TensorLoad.scala 202:86:@2974.6]
  reg [9:0] waddr_cur; // @[TensorLoad.scala 206:22:@2979.4]
  reg [31:0] _RAND_36;
  reg [9:0] waddr_nxt; // @[TensorLoad.scala 207:22:@2980.4]
  reg [31:0] _RAND_37;
  wire  _T_4523; // @[TensorLoad.scala 212:5:@2990.6]
  wire  _T_4526; // @[TensorLoad.scala 213:5:@2992.6]
  wire [10:0] _T_4528; // @[TensorLoad.scala 215:28:@2994.8]
  wire [9:0] _T_4529; // @[TensorLoad.scala 215:28:@2995.8]
  wire  _T_4531; // @[TensorLoad.scala 216:33:@3000.8]
  wire [15:0] _GEN_426; // @[TensorLoad.scala 217:28:@3002.10]
  wire [16:0] _T_4532; // @[TensorLoad.scala 217:28:@3002.10]
  wire [15:0] _T_4533; // @[TensorLoad.scala 217:28:@3003.10]
  wire [15:0] _GEN_33; // @[TensorLoad.scala 216:59:@3001.8]
  wire [15:0] _GEN_34; // @[TensorLoad.scala 216:59:@3001.8]
  wire [15:0] _GEN_35; // @[TensorLoad.scala 214:3:@2993.6]
  wire [15:0] _GEN_36; // @[TensorLoad.scala 214:3:@2993.6]
  wire [15:0] _GEN_37; // @[TensorLoad.scala 208:25:@2982.4]
  wire [15:0] _GEN_38; // @[TensorLoad.scala 208:25:@2982.4]
  wire  wmask_0_0; // @[TensorLoad.scala 235:26:@3060.4]
  wire [63:0] wdata_0_0; // @[TensorLoad.scala 236:25:@3062.4]
  wire  _T_4947; // @[TensorLoad.scala 242:51:@3093.4]
  wire  _T_4948; // @[TensorLoad.scala 242:45:@3094.4]
  wire  _T_5034; // @[TensorLoad.scala 242:51:@3144.4]
  wire  _T_5035; // @[TensorLoad.scala 242:45:@3145.4]
  wire  _T_5121; // @[TensorLoad.scala 242:51:@3195.4]
  wire  _T_5122; // @[TensorLoad.scala 242:45:@3196.4]
  wire  _T_5208; // @[TensorLoad.scala 242:51:@3246.4]
  wire  _T_5209; // @[TensorLoad.scala 242:45:@3247.4]
  wire  _T_5295; // @[TensorLoad.scala 242:51:@3297.4]
  wire  _T_5296; // @[TensorLoad.scala 242:45:@3298.4]
  wire  _T_5382; // @[TensorLoad.scala 242:51:@3348.4]
  wire  _T_5383; // @[TensorLoad.scala 242:45:@3349.4]
  wire  _T_5469; // @[TensorLoad.scala 242:51:@3399.4]
  wire  _T_5470; // @[TensorLoad.scala 242:45:@3400.4]
  wire  _T_5556; // @[TensorLoad.scala 242:51:@3450.4]
  wire  _T_5557; // @[TensorLoad.scala 242:45:@3451.4]
  wire  _T_5643; // @[TensorLoad.scala 242:51:@3501.4]
  wire  _T_5644; // @[TensorLoad.scala 242:45:@3502.4]
  wire  _T_5730; // @[TensorLoad.scala 242:51:@3552.4]
  wire  _T_5731; // @[TensorLoad.scala 242:45:@3553.4]
  wire  _T_5817; // @[TensorLoad.scala 242:51:@3603.4]
  wire  _T_5818; // @[TensorLoad.scala 242:45:@3604.4]
  wire  _T_5904; // @[TensorLoad.scala 242:51:@3654.4]
  wire  _T_5905; // @[TensorLoad.scala 242:45:@3655.4]
  wire  _T_5991; // @[TensorLoad.scala 242:51:@3705.4]
  wire  _T_5992; // @[TensorLoad.scala 242:45:@3706.4]
  wire  _T_6078; // @[TensorLoad.scala 242:51:@3756.4]
  wire  _T_6079; // @[TensorLoad.scala 242:45:@3757.4]
  wire  _T_6165; // @[TensorLoad.scala 242:51:@3807.4]
  wire  _T_6166; // @[TensorLoad.scala 242:45:@3808.4]
  reg  rvalid; // @[TensorLoad.scala 252:23:@3876.4]
  reg [31:0] _RAND_38;
  wire  _GEN_216; // @[TensorLoad.scala 256:26:@3881.4]
  wire [127:0] _T_6482; // @[TensorLoad.scala 259:38:@4007.4]
  wire [127:0] _T_6624; // @[TensorLoad.scala 259:38:@4059.4]
  wire [127:0] _T_6766; // @[TensorLoad.scala 259:38:@4111.4]
  wire [127:0] _T_6908; // @[TensorLoad.scala 259:38:@4163.4]
  wire [127:0] _T_7050; // @[TensorLoad.scala 259:38:@4215.4]
  wire [127:0] _T_7192; // @[TensorLoad.scala 259:38:@4267.4]
  wire [127:0] _T_7334; // @[TensorLoad.scala 259:38:@4319.4]
  wire [127:0] _T_7476; // @[TensorLoad.scala 259:38:@4371.4]
  wire [127:0] _T_7618; // @[TensorLoad.scala 259:38:@4423.4]
  wire [127:0] _T_7760; // @[TensorLoad.scala 259:38:@4475.4]
  wire [127:0] _T_7902; // @[TensorLoad.scala 259:38:@4527.4]
  wire [127:0] _T_8044; // @[TensorLoad.scala 259:38:@4579.4]
  wire [127:0] _T_8186; // @[TensorLoad.scala 259:38:@4631.4]
  wire [127:0] _T_8328; // @[TensorLoad.scala 259:38:@4683.4]
  wire [127:0] _T_8470; // @[TensorLoad.scala 259:38:@4735.4]
  wire [127:0] _T_8612; // @[TensorLoad.scala 259:38:@4787.4]
  wire  _T_8760; // @[TensorLoad.scala 263:96:@4843.4]
  wire  done_no_pad; // @[TensorLoad.scala 263:83:@4844.4]
  wire  done_x_pad; // @[TensorLoad.scala 264:72:@4849.4]
  wire  _T_8767; // @[TensorLoad.scala 265:37:@4851.4]
  wire  done_y_pad; // @[TensorLoad.scala 265:52:@4852.4]
  wire  _T_8768; // @[TensorLoad.scala 266:26:@4853.4]
  reg [9:0] tensorFile_0_0_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_39;
  reg [9:0] tensorFile_0_1_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_40;
  reg [9:0] tensorFile_1_0_rdata_1_addr_pipe_0;
  reg [31:0] _RAND_41;
  reg [9:0] tensorFile_1_1_rdata_1_addr_pipe_0;
  reg [31:0] _RAND_42;
  reg [9:0] tensorFile_2_0_rdata_2_addr_pipe_0;
  reg [31:0] _RAND_43;
  reg [9:0] tensorFile_2_1_rdata_2_addr_pipe_0;
  reg [31:0] _RAND_44;
  reg [9:0] tensorFile_3_0_rdata_3_addr_pipe_0;
  reg [31:0] _RAND_45;
  reg [9:0] tensorFile_3_1_rdata_3_addr_pipe_0;
  reg [31:0] _RAND_46;
  reg [9:0] tensorFile_4_0_rdata_4_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [9:0] tensorFile_4_1_rdata_4_addr_pipe_0;
  reg [31:0] _RAND_48;
  reg [9:0] tensorFile_5_0_rdata_5_addr_pipe_0;
  reg [31:0] _RAND_49;
  reg [9:0] tensorFile_5_1_rdata_5_addr_pipe_0;
  reg [31:0] _RAND_50;
  reg [9:0] tensorFile_6_0_rdata_6_addr_pipe_0;
  reg [31:0] _RAND_51;
  reg [9:0] tensorFile_6_1_rdata_6_addr_pipe_0;
  reg [31:0] _RAND_52;
  reg [9:0] tensorFile_7_0_rdata_7_addr_pipe_0;
  reg [31:0] _RAND_53;
  reg [9:0] tensorFile_7_1_rdata_7_addr_pipe_0;
  reg [31:0] _RAND_54;
  reg [9:0] tensorFile_8_0_rdata_8_addr_pipe_0;
  reg [31:0] _RAND_55;
  reg [9:0] tensorFile_8_1_rdata_8_addr_pipe_0;
  reg [31:0] _RAND_56;
  reg [9:0] tensorFile_9_0_rdata_9_addr_pipe_0;
  reg [31:0] _RAND_57;
  reg [9:0] tensorFile_9_1_rdata_9_addr_pipe_0;
  reg [31:0] _RAND_58;
  reg [9:0] tensorFile_10_0_rdata_10_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [9:0] tensorFile_10_1_rdata_10_addr_pipe_0;
  reg [31:0] _RAND_60;
  reg [9:0] tensorFile_11_0_rdata_11_addr_pipe_0;
  reg [31:0] _RAND_61;
  reg [9:0] tensorFile_11_1_rdata_11_addr_pipe_0;
  reg [31:0] _RAND_62;
  reg [9:0] tensorFile_12_0_rdata_12_addr_pipe_0;
  reg [31:0] _RAND_63;
  reg [9:0] tensorFile_12_1_rdata_12_addr_pipe_0;
  reg [31:0] _RAND_64;
  reg [9:0] tensorFile_13_0_rdata_13_addr_pipe_0;
  reg [31:0] _RAND_65;
  reg [9:0] tensorFile_13_1_rdata_13_addr_pipe_0;
  reg [31:0] _RAND_66;
  reg [9:0] tensorFile_14_0_rdata_14_addr_pipe_0;
  reg [31:0] _RAND_67;
  reg [9:0] tensorFile_14_1_rdata_14_addr_pipe_0;
  reg [31:0] _RAND_68;
  reg [9:0] tensorFile_15_0_rdata_15_addr_pipe_0;
  reg [31:0] _RAND_69;
  reg [9:0] tensorFile_15_1_rdata_15_addr_pipe_0;
  reg [31:0] _RAND_70;
  TensorDataCtrl_1 dataCtrl ( // @[TensorLoad.scala 52:24:@2726.4]
    .clock(dataCtrl_clock),
    .io_start(dataCtrl_io_start),
    .io_done(dataCtrl_io_done),
    .io_inst(dataCtrl_io_inst),
    .io_baddr(dataCtrl_io_baddr),
    .io_xinit(dataCtrl_io_xinit),
    .io_xupdate(dataCtrl_io_xupdate),
    .io_yupdate(dataCtrl_io_yupdate),
    .io_stride(dataCtrl_io_stride),
    .io_split(dataCtrl_io_split),
    .io_addr(dataCtrl_io_addr),
    .io_len(dataCtrl_io_len)
  );
  TensorPadCtrl_4 yPadCtrl0 ( // @[TensorLoad.scala 55:25:@2730.4]
    .clock(yPadCtrl0_clock),
    .reset(yPadCtrl0_reset),
    .io_start(yPadCtrl0_io_start),
    .io_done(yPadCtrl0_io_done),
    .io_inst(yPadCtrl0_io_inst)
  );
  TensorPadCtrl_5 yPadCtrl1 ( // @[TensorLoad.scala 56:25:@2733.4]
    .clock(yPadCtrl1_clock),
    .reset(yPadCtrl1_reset),
    .io_start(yPadCtrl1_io_start),
    .io_done(yPadCtrl1_io_done),
    .io_inst(yPadCtrl1_io_inst)
  );
  TensorPadCtrl_6 xPadCtrl0 ( // @[TensorLoad.scala 57:25:@2736.4]
    .clock(xPadCtrl0_clock),
    .reset(xPadCtrl0_reset),
    .io_start(xPadCtrl0_io_start),
    .io_done(xPadCtrl0_io_done),
    .io_inst(xPadCtrl0_io_inst)
  );
  TensorPadCtrl_7 xPadCtrl1 ( // @[TensorLoad.scala 58:25:@2739.4]
    .clock(xPadCtrl1_clock),
    .reset(xPadCtrl1_reset),
    .io_start(xPadCtrl1_io_start),
    .io_done(xPadCtrl1_io_done),
    .io_inst(xPadCtrl1_io_inst)
  );
  assign tensorFile_0_0_rdata_0_addr = tensorFile_0_0_rdata_0_addr_pipe_0;
  assign tensorFile_0_0_rdata_0_data = tensorFile_0_0[tensorFile_0_0_rdata_0_addr]; // @[TensorLoad.scala 222:16:@3009.4]
  assign tensorFile_0_0__T_4976_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_0_0__T_4976_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_0_0__T_4976_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_0_0__T_4976_en = _T_4420 ? 1'h0 : _T_4948;
  assign tensorFile_0_1_rdata_0_addr = tensorFile_0_1_rdata_0_addr_pipe_0;
  assign tensorFile_0_1_rdata_0_data = tensorFile_0_1[tensorFile_0_1_rdata_0_addr]; // @[TensorLoad.scala 222:16:@3009.4]
  assign tensorFile_0_1__T_4976_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_0_1__T_4976_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_0_1__T_4976_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_0_1__T_4976_en = _T_4420 ? 1'h0 : _T_4948;
  assign tensorFile_1_0_rdata_1_addr = tensorFile_1_0_rdata_1_addr_pipe_0;
  assign tensorFile_1_0_rdata_1_data = tensorFile_1_0[tensorFile_1_0_rdata_1_addr]; // @[TensorLoad.scala 222:16:@3010.4]
  assign tensorFile_1_0__T_5063_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_1_0__T_5063_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_1_0__T_5063_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_1_0__T_5063_en = _T_4420 ? 1'h0 : _T_5035;
  assign tensorFile_1_1_rdata_1_addr = tensorFile_1_1_rdata_1_addr_pipe_0;
  assign tensorFile_1_1_rdata_1_data = tensorFile_1_1[tensorFile_1_1_rdata_1_addr]; // @[TensorLoad.scala 222:16:@3010.4]
  assign tensorFile_1_1__T_5063_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_1_1__T_5063_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_1_1__T_5063_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_1_1__T_5063_en = _T_4420 ? 1'h0 : _T_5035;
  assign tensorFile_2_0_rdata_2_addr = tensorFile_2_0_rdata_2_addr_pipe_0;
  assign tensorFile_2_0_rdata_2_data = tensorFile_2_0[tensorFile_2_0_rdata_2_addr]; // @[TensorLoad.scala 222:16:@3011.4]
  assign tensorFile_2_0__T_5150_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_2_0__T_5150_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_2_0__T_5150_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_2_0__T_5150_en = _T_4420 ? 1'h0 : _T_5122;
  assign tensorFile_2_1_rdata_2_addr = tensorFile_2_1_rdata_2_addr_pipe_0;
  assign tensorFile_2_1_rdata_2_data = tensorFile_2_1[tensorFile_2_1_rdata_2_addr]; // @[TensorLoad.scala 222:16:@3011.4]
  assign tensorFile_2_1__T_5150_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_2_1__T_5150_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_2_1__T_5150_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_2_1__T_5150_en = _T_4420 ? 1'h0 : _T_5122;
  assign tensorFile_3_0_rdata_3_addr = tensorFile_3_0_rdata_3_addr_pipe_0;
  assign tensorFile_3_0_rdata_3_data = tensorFile_3_0[tensorFile_3_0_rdata_3_addr]; // @[TensorLoad.scala 222:16:@3012.4]
  assign tensorFile_3_0__T_5237_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_3_0__T_5237_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_3_0__T_5237_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_3_0__T_5237_en = _T_4420 ? 1'h0 : _T_5209;
  assign tensorFile_3_1_rdata_3_addr = tensorFile_3_1_rdata_3_addr_pipe_0;
  assign tensorFile_3_1_rdata_3_data = tensorFile_3_1[tensorFile_3_1_rdata_3_addr]; // @[TensorLoad.scala 222:16:@3012.4]
  assign tensorFile_3_1__T_5237_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_3_1__T_5237_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_3_1__T_5237_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_3_1__T_5237_en = _T_4420 ? 1'h0 : _T_5209;
  assign tensorFile_4_0_rdata_4_addr = tensorFile_4_0_rdata_4_addr_pipe_0;
  assign tensorFile_4_0_rdata_4_data = tensorFile_4_0[tensorFile_4_0_rdata_4_addr]; // @[TensorLoad.scala 222:16:@3013.4]
  assign tensorFile_4_0__T_5324_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_4_0__T_5324_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_4_0__T_5324_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_4_0__T_5324_en = _T_4420 ? 1'h0 : _T_5296;
  assign tensorFile_4_1_rdata_4_addr = tensorFile_4_1_rdata_4_addr_pipe_0;
  assign tensorFile_4_1_rdata_4_data = tensorFile_4_1[tensorFile_4_1_rdata_4_addr]; // @[TensorLoad.scala 222:16:@3013.4]
  assign tensorFile_4_1__T_5324_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_4_1__T_5324_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_4_1__T_5324_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_4_1__T_5324_en = _T_4420 ? 1'h0 : _T_5296;
  assign tensorFile_5_0_rdata_5_addr = tensorFile_5_0_rdata_5_addr_pipe_0;
  assign tensorFile_5_0_rdata_5_data = tensorFile_5_0[tensorFile_5_0_rdata_5_addr]; // @[TensorLoad.scala 222:16:@3014.4]
  assign tensorFile_5_0__T_5411_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_5_0__T_5411_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_5_0__T_5411_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_5_0__T_5411_en = _T_4420 ? 1'h0 : _T_5383;
  assign tensorFile_5_1_rdata_5_addr = tensorFile_5_1_rdata_5_addr_pipe_0;
  assign tensorFile_5_1_rdata_5_data = tensorFile_5_1[tensorFile_5_1_rdata_5_addr]; // @[TensorLoad.scala 222:16:@3014.4]
  assign tensorFile_5_1__T_5411_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_5_1__T_5411_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_5_1__T_5411_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_5_1__T_5411_en = _T_4420 ? 1'h0 : _T_5383;
  assign tensorFile_6_0_rdata_6_addr = tensorFile_6_0_rdata_6_addr_pipe_0;
  assign tensorFile_6_0_rdata_6_data = tensorFile_6_0[tensorFile_6_0_rdata_6_addr]; // @[TensorLoad.scala 222:16:@3015.4]
  assign tensorFile_6_0__T_5498_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_6_0__T_5498_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_6_0__T_5498_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_6_0__T_5498_en = _T_4420 ? 1'h0 : _T_5470;
  assign tensorFile_6_1_rdata_6_addr = tensorFile_6_1_rdata_6_addr_pipe_0;
  assign tensorFile_6_1_rdata_6_data = tensorFile_6_1[tensorFile_6_1_rdata_6_addr]; // @[TensorLoad.scala 222:16:@3015.4]
  assign tensorFile_6_1__T_5498_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_6_1__T_5498_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_6_1__T_5498_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_6_1__T_5498_en = _T_4420 ? 1'h0 : _T_5470;
  assign tensorFile_7_0_rdata_7_addr = tensorFile_7_0_rdata_7_addr_pipe_0;
  assign tensorFile_7_0_rdata_7_data = tensorFile_7_0[tensorFile_7_0_rdata_7_addr]; // @[TensorLoad.scala 222:16:@3016.4]
  assign tensorFile_7_0__T_5585_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_7_0__T_5585_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_7_0__T_5585_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_7_0__T_5585_en = _T_4420 ? 1'h0 : _T_5557;
  assign tensorFile_7_1_rdata_7_addr = tensorFile_7_1_rdata_7_addr_pipe_0;
  assign tensorFile_7_1_rdata_7_data = tensorFile_7_1[tensorFile_7_1_rdata_7_addr]; // @[TensorLoad.scala 222:16:@3016.4]
  assign tensorFile_7_1__T_5585_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_7_1__T_5585_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_7_1__T_5585_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_7_1__T_5585_en = _T_4420 ? 1'h0 : _T_5557;
  assign tensorFile_8_0_rdata_8_addr = tensorFile_8_0_rdata_8_addr_pipe_0;
  assign tensorFile_8_0_rdata_8_data = tensorFile_8_0[tensorFile_8_0_rdata_8_addr]; // @[TensorLoad.scala 222:16:@3017.4]
  assign tensorFile_8_0__T_5672_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_8_0__T_5672_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_8_0__T_5672_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_8_0__T_5672_en = _T_4420 ? 1'h0 : _T_5644;
  assign tensorFile_8_1_rdata_8_addr = tensorFile_8_1_rdata_8_addr_pipe_0;
  assign tensorFile_8_1_rdata_8_data = tensorFile_8_1[tensorFile_8_1_rdata_8_addr]; // @[TensorLoad.scala 222:16:@3017.4]
  assign tensorFile_8_1__T_5672_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_8_1__T_5672_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_8_1__T_5672_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_8_1__T_5672_en = _T_4420 ? 1'h0 : _T_5644;
  assign tensorFile_9_0_rdata_9_addr = tensorFile_9_0_rdata_9_addr_pipe_0;
  assign tensorFile_9_0_rdata_9_data = tensorFile_9_0[tensorFile_9_0_rdata_9_addr]; // @[TensorLoad.scala 222:16:@3018.4]
  assign tensorFile_9_0__T_5759_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_9_0__T_5759_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_9_0__T_5759_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_9_0__T_5759_en = _T_4420 ? 1'h0 : _T_5731;
  assign tensorFile_9_1_rdata_9_addr = tensorFile_9_1_rdata_9_addr_pipe_0;
  assign tensorFile_9_1_rdata_9_data = tensorFile_9_1[tensorFile_9_1_rdata_9_addr]; // @[TensorLoad.scala 222:16:@3018.4]
  assign tensorFile_9_1__T_5759_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_9_1__T_5759_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_9_1__T_5759_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_9_1__T_5759_en = _T_4420 ? 1'h0 : _T_5731;
  assign tensorFile_10_0_rdata_10_addr = tensorFile_10_0_rdata_10_addr_pipe_0;
  assign tensorFile_10_0_rdata_10_data = tensorFile_10_0[tensorFile_10_0_rdata_10_addr]; // @[TensorLoad.scala 222:16:@3019.4]
  assign tensorFile_10_0__T_5846_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_10_0__T_5846_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_10_0__T_5846_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_10_0__T_5846_en = _T_4420 ? 1'h0 : _T_5818;
  assign tensorFile_10_1_rdata_10_addr = tensorFile_10_1_rdata_10_addr_pipe_0;
  assign tensorFile_10_1_rdata_10_data = tensorFile_10_1[tensorFile_10_1_rdata_10_addr]; // @[TensorLoad.scala 222:16:@3019.4]
  assign tensorFile_10_1__T_5846_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_10_1__T_5846_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_10_1__T_5846_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_10_1__T_5846_en = _T_4420 ? 1'h0 : _T_5818;
  assign tensorFile_11_0_rdata_11_addr = tensorFile_11_0_rdata_11_addr_pipe_0;
  assign tensorFile_11_0_rdata_11_data = tensorFile_11_0[tensorFile_11_0_rdata_11_addr]; // @[TensorLoad.scala 222:16:@3020.4]
  assign tensorFile_11_0__T_5933_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_11_0__T_5933_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_11_0__T_5933_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_11_0__T_5933_en = _T_4420 ? 1'h0 : _T_5905;
  assign tensorFile_11_1_rdata_11_addr = tensorFile_11_1_rdata_11_addr_pipe_0;
  assign tensorFile_11_1_rdata_11_data = tensorFile_11_1[tensorFile_11_1_rdata_11_addr]; // @[TensorLoad.scala 222:16:@3020.4]
  assign tensorFile_11_1__T_5933_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_11_1__T_5933_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_11_1__T_5933_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_11_1__T_5933_en = _T_4420 ? 1'h0 : _T_5905;
  assign tensorFile_12_0_rdata_12_addr = tensorFile_12_0_rdata_12_addr_pipe_0;
  assign tensorFile_12_0_rdata_12_data = tensorFile_12_0[tensorFile_12_0_rdata_12_addr]; // @[TensorLoad.scala 222:16:@3021.4]
  assign tensorFile_12_0__T_6020_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_12_0__T_6020_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_12_0__T_6020_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_12_0__T_6020_en = _T_4420 ? 1'h0 : _T_5992;
  assign tensorFile_12_1_rdata_12_addr = tensorFile_12_1_rdata_12_addr_pipe_0;
  assign tensorFile_12_1_rdata_12_data = tensorFile_12_1[tensorFile_12_1_rdata_12_addr]; // @[TensorLoad.scala 222:16:@3021.4]
  assign tensorFile_12_1__T_6020_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_12_1__T_6020_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_12_1__T_6020_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_12_1__T_6020_en = _T_4420 ? 1'h0 : _T_5992;
  assign tensorFile_13_0_rdata_13_addr = tensorFile_13_0_rdata_13_addr_pipe_0;
  assign tensorFile_13_0_rdata_13_data = tensorFile_13_0[tensorFile_13_0_rdata_13_addr]; // @[TensorLoad.scala 222:16:@3022.4]
  assign tensorFile_13_0__T_6107_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_13_0__T_6107_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_13_0__T_6107_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_13_0__T_6107_en = _T_4420 ? 1'h0 : _T_6079;
  assign tensorFile_13_1_rdata_13_addr = tensorFile_13_1_rdata_13_addr_pipe_0;
  assign tensorFile_13_1_rdata_13_data = tensorFile_13_1[tensorFile_13_1_rdata_13_addr]; // @[TensorLoad.scala 222:16:@3022.4]
  assign tensorFile_13_1__T_6107_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_13_1__T_6107_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_13_1__T_6107_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_13_1__T_6107_en = _T_4420 ? 1'h0 : _T_6079;
  assign tensorFile_14_0_rdata_14_addr = tensorFile_14_0_rdata_14_addr_pipe_0;
  assign tensorFile_14_0_rdata_14_data = tensorFile_14_0[tensorFile_14_0_rdata_14_addr]; // @[TensorLoad.scala 222:16:@3023.4]
  assign tensorFile_14_0__T_6194_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_14_0__T_6194_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_14_0__T_6194_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_14_0__T_6194_en = _T_4420 ? 1'h0 : _T_6166;
  assign tensorFile_14_1_rdata_14_addr = tensorFile_14_1_rdata_14_addr_pipe_0;
  assign tensorFile_14_1_rdata_14_data = tensorFile_14_1[tensorFile_14_1_rdata_14_addr]; // @[TensorLoad.scala 222:16:@3023.4]
  assign tensorFile_14_1__T_6194_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_14_1__T_6194_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_14_1__T_6194_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_14_1__T_6194_en = _T_4420 ? 1'h0 : _T_6166;
  assign tensorFile_15_0_rdata_15_addr = tensorFile_15_0_rdata_15_addr_pipe_0;
  assign tensorFile_15_0_rdata_15_data = tensorFile_15_0[tensorFile_15_0_rdata_15_addr]; // @[TensorLoad.scala 222:16:@3024.4]
  assign tensorFile_15_0__T_6281_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_15_0__T_6281_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_15_0__T_6281_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_15_0__T_6281_en = _T_4420 ? 1'h0 : _T_4523;
  assign tensorFile_15_1_rdata_15_addr = tensorFile_15_1_rdata_15_addr_pipe_0;
  assign tensorFile_15_1_rdata_15_data = tensorFile_15_1[tensorFile_15_1_rdata_15_addr]; // @[TensorLoad.scala 222:16:@3024.4]
  assign tensorFile_15_1__T_6281_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_15_1__T_6281_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_15_1__T_6281_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_15_1__T_6281_en = _T_4420 ? 1'h0 : _T_4523;
  assign dec_sram_offset = io_inst[24:9]; // @[TensorLoad.scala 51:29:@2706.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorLoad.scala 51:29:@2714.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorLoad.scala 51:29:@2718.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorLoad.scala 51:29:@2720.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorLoad.scala 51:29:@2722.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorLoad.scala 51:29:@2724.4]
  assign _T_4394 = 3'h0 == state; // @[Conditional.scala 37:30:@2745.4]
  assign _T_4396 = dec_ypad_0 != 4'h0; // @[TensorLoad.scala 71:25:@2748.8]
  assign _T_4398 = dec_xpad_0 != 4'h0; // @[TensorLoad.scala 73:31:@2753.10]
  assign _GEN_0 = _T_4398 ? 3'h2 : 3'h3; // @[TensorLoad.scala 73:40:@2754.10]
  assign _GEN_1 = _T_4396 ? 3'h1 : _GEN_0; // @[TensorLoad.scala 71:34:@2749.8]
  assign _GEN_2 = io_start ? _GEN_1 : state; // @[TensorLoad.scala 70:22:@2747.6]
  assign _T_4399 = 3'h1 == state; // @[Conditional.scala 37:30:@2763.6]
  assign _GEN_4 = yPadCtrl0_io_done ? _GEN_0 : state; // @[TensorLoad.scala 81:31:@2765.8]
  assign _T_4402 = 3'h2 == state; // @[Conditional.scala 37:30:@2776.8]
  assign _GEN_5 = xPadCtrl0_io_done ? 3'h3 : state; // @[TensorLoad.scala 90:31:@2778.10]
  assign _T_4403 = 3'h3 == state; // @[Conditional.scala 37:30:@2783.10]
  assign _GEN_6 = io_vme_rd_cmd_ready ? 3'h4 : state; // @[TensorLoad.scala 95:33:@2785.12]
  assign _T_4404 = 3'h4 == state; // @[Conditional.scala 37:30:@2790.12]
  assign _T_4406 = dec_xpad_1 != 4'h0; // @[TensorLoad.scala 102:27:@2794.18]
  assign _T_4408 = dec_ypad_1 != 4'h0; // @[TensorLoad.scala 104:33:@2799.20]
  assign _GEN_7 = _T_4408 ? 3'h6 : 3'h0; // @[TensorLoad.scala 104:42:@2800.20]
  assign _GEN_8 = _T_4406 ? 3'h5 : _GEN_7; // @[TensorLoad.scala 102:36:@2795.18]
  assign _GEN_10 = _T_4406 ? 3'h5 : _GEN_0; // @[TensorLoad.scala 110:36:@2810.20]
  assign _GEN_11 = dataCtrl_io_split ? 3'h3 : state; // @[TensorLoad.scala 117:39:@2823.20]
  assign _GEN_12 = dataCtrl_io_stride ? _GEN_10 : _GEN_11; // @[TensorLoad.scala 109:40:@2808.18]
  assign _GEN_13 = dataCtrl_io_done ? _GEN_8 : _GEN_12; // @[TensorLoad.scala 101:32:@2793.16]
  assign _GEN_14 = io_vme_rd_data_valid ? _GEN_13 : state; // @[TensorLoad.scala 100:34:@2792.14]
  assign _T_4413 = 3'h5 == state; // @[Conditional.scala 37:30:@2829.14]
  assign _GEN_17 = dataCtrlDone ? _GEN_7 : _GEN_0; // @[TensorLoad.scala 124:28:@2832.18]
  assign _GEN_18 = xPadCtrl1_io_done ? _GEN_17 : state; // @[TensorLoad.scala 123:31:@2831.16]
  assign _T_4418 = 3'h6 == state; // @[Conditional.scala 37:30:@2853.16]
  assign _T_4419 = yPadCtrl1_io_done & dataCtrlDone; // @[TensorLoad.scala 140:30:@2855.18]
  assign _GEN_19 = _T_4419 ? 3'h0 : state; // @[TensorLoad.scala 140:47:@2856.18]
  assign _GEN_20 = _T_4418 ? _GEN_19 : state; // @[Conditional.scala 39:67:@2854.16]
  assign _GEN_21 = _T_4413 ? _GEN_18 : _GEN_20; // @[Conditional.scala 39:67:@2830.14]
  assign _GEN_22 = _T_4404 ? _GEN_14 : _GEN_21; // @[Conditional.scala 39:67:@2791.12]
  assign _GEN_23 = _T_4403 ? _GEN_6 : _GEN_22; // @[Conditional.scala 39:67:@2784.10]
  assign _GEN_24 = _T_4402 ? _GEN_5 : _GEN_23; // @[Conditional.scala 39:67:@2777.8]
  assign _GEN_25 = _T_4399 ? _GEN_4 : _GEN_24; // @[Conditional.scala 39:67:@2764.6]
  assign _GEN_26 = _T_4394 ? _GEN_2 : _GEN_25; // @[Conditional.scala 40:58:@2746.4]
  assign _T_4420 = state == 3'h0; // @[TensorLoad.scala 147:30:@2860.4]
  assign _T_4421 = _T_4420 & io_start; // @[TensorLoad.scala 147:40:@2861.4]
  assign _T_4423 = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[Decoupled.scala 37:37:@2867.4]
  assign _T_4428 = _T_4423 & dataCtrl_io_done; // @[TensorLoad.scala 156:36:@2877.6]
  assign _GEN_27 = _T_4428 ? 1'h1 : dataCtrlDone; // @[TensorLoad.scala 156:57:@2878.6]
  assign _GEN_28 = _T_4420 ? 1'h0 : _GEN_27; // @[TensorLoad.scala 154:25:@2872.4]
  assign _T_4433 = _T_4396 & _T_4420; // @[TensorLoad.scala 161:44:@2883.4]
  assign _T_4440 = dec_xpad_1 == 4'h0; // @[TensorLoad.scala 164:61:@2889.4]
  assign _T_4441 = _T_4428 & _T_4440; // @[TensorLoad.scala 164:48:@2890.4]
  assign _T_4442 = state == 3'h5; // @[TensorLoad.scala 165:14:@2891.4]
  assign _T_4443 = _T_4442 & xPadCtrl1_io_done; // @[TensorLoad.scala 165:25:@2892.4]
  assign _T_4444 = _T_4443 & dataCtrlDone; // @[TensorLoad.scala 165:45:@2893.4]
  assign _T_4445 = _T_4441 | _T_4444; // @[TensorLoad.scala 164:70:@2894.4]
  assign _T_4451 = state == 3'h1; // @[TensorLoad.scala 169:14:@2900.4]
  assign _T_4452 = _T_4451 & yPadCtrl0_io_done; // @[TensorLoad.scala 169:25:@2901.4]
  assign _T_4453 = _T_4421 | _T_4452; // @[TensorLoad.scala 168:35:@2902.4]
  assign _T_4455 = ~ dataCtrlDone; // @[TensorLoad.scala 170:32:@2904.4]
  assign _T_4456 = _T_4423 & _T_4455; // @[TensorLoad.scala 170:30:@2905.4]
  assign _T_4457 = _T_4456 & dataCtrl_io_stride; // @[TensorLoad.scala 170:46:@2906.4]
  assign _T_4460 = _T_4457 & _T_4440; // @[TensorLoad.scala 170:67:@2908.4]
  assign _T_4461 = _T_4453 | _T_4460; // @[TensorLoad.scala 169:46:@2909.4]
  assign _T_4465 = _T_4443 & _T_4455; // @[TensorLoad.scala 171:45:@2913.4]
  assign _T_4466 = _T_4461 | _T_4465; // @[TensorLoad.scala 170:89:@2914.4]
  assign _T_4471 = _T_4406 & _T_4423; // @[TensorLoad.scala 173:44:@2919.4]
  assign _T_4472 = ~ dataCtrl_io_done; // @[TensorLoad.scala 174:28:@2920.4]
  assign _T_4473 = _T_4472 & dataCtrl_io_stride; // @[TensorLoad.scala 174:46:@2921.4]
  assign _T_4476 = _T_4473 & _T_4406; // @[TensorLoad.scala 174:67:@2923.4]
  assign _T_4477 = dataCtrl_io_done | _T_4476; // @[TensorLoad.scala 174:25:@2924.4]
  assign _T_4479 = state == 3'h3; // @[TensorLoad.scala 182:32:@2931.4]
  assign _T_4482 = state == 3'h2; // @[TensorLoad.scala 190:11:@2938.4]
  assign _T_4483 = _T_4451 | _T_4482; // @[TensorLoad.scala 189:36:@2939.4]
  assign _T_4485 = _T_4483 | _T_4442; // @[TensorLoad.scala 190:22:@2941.4]
  assign _T_4486 = state == 3'h6; // @[TensorLoad.scala 192:11:@2942.4]
  assign isZeroPad = _T_4485 | _T_4486; // @[TensorLoad.scala 191:22:@2943.4]
  assign _T_4489 = _T_4420 | _T_4479; // @[TensorLoad.scala 194:24:@2946.4]
  assign _T_4492 = _T_4489 | tag; // @[TensorLoad.scala 194:46:@2948.4]
  assign _T_4495 = _T_4423 | isZeroPad; // @[TensorLoad.scala 196:36:@2954.6]
  assign _T_4497 = tag + 1'h1; // @[TensorLoad.scala 197:16:@2956.8]
  assign _T_4498 = tag + 1'h1; // @[TensorLoad.scala 197:16:@2957.8]
  assign _GEN_29 = _T_4495 ? _T_4498 : tag; // @[TensorLoad.scala 196:50:@2955.6]
  assign _T_4500 = _T_4420 | dataCtrlDone; // @[TensorLoad.scala 200:24:@2961.4]
  assign _T_4502 = set == 4'hf; // @[TensorLoad.scala 200:48:@2962.4]
  assign _T_4505 = _T_4502 & tag; // @[TensorLoad.scala 200:76:@2964.4]
  assign _T_4506 = _T_4500 | _T_4505; // @[TensorLoad.scala 200:40:@2965.4]
  assign _T_4512 = _T_4495 & tag; // @[TensorLoad.scala 202:51:@2973.6]
  assign _T_4514 = set + 4'h1; // @[TensorLoad.scala 203:16:@2975.8]
  assign _T_4515 = set + 4'h1; // @[TensorLoad.scala 203:16:@2976.8]
  assign _GEN_31 = _T_4512 ? _T_4515 : set; // @[TensorLoad.scala 202:86:@2974.6]
  assign _T_4523 = _T_4495 & _T_4502; // @[TensorLoad.scala 212:5:@2990.6]
  assign _T_4526 = _T_4523 & tag; // @[TensorLoad.scala 213:5:@2992.6]
  assign _T_4528 = waddr_cur + 10'h1; // @[TensorLoad.scala 215:28:@2994.8]
  assign _T_4529 = waddr_cur + 10'h1; // @[TensorLoad.scala 215:28:@2995.8]
  assign _T_4531 = dataCtrl_io_stride & _T_4423; // @[TensorLoad.scala 216:33:@3000.8]
  assign _GEN_426 = {{6'd0}, waddr_nxt}; // @[TensorLoad.scala 217:28:@3002.10]
  assign _T_4532 = _GEN_426 + dec_xsize; // @[TensorLoad.scala 217:28:@3002.10]
  assign _T_4533 = _GEN_426 + dec_xsize; // @[TensorLoad.scala 217:28:@3003.10]
  assign _GEN_33 = _T_4531 ? _T_4533 : {{6'd0}, waddr_cur}; // @[TensorLoad.scala 216:59:@3001.8]
  assign _GEN_34 = _T_4531 ? _T_4533 : {{6'd0}, waddr_nxt}; // @[TensorLoad.scala 216:59:@3001.8]
  assign _GEN_35 = _T_4526 ? {{6'd0}, _T_4529} : _GEN_33; // @[TensorLoad.scala 214:3:@2993.6]
  assign _GEN_36 = _T_4526 ? {{6'd0}, waddr_nxt} : _GEN_34; // @[TensorLoad.scala 214:3:@2993.6]
  assign _GEN_37 = _T_4420 ? dec_sram_offset : _GEN_35; // @[TensorLoad.scala 208:25:@2982.4]
  assign _GEN_38 = _T_4420 ? dec_sram_offset : _GEN_36; // @[TensorLoad.scala 208:25:@2982.4]
  assign wmask_0_0 = tag == 1'h0; // @[TensorLoad.scala 235:26:@3060.4]
  assign wdata_0_0 = isZeroPad ? 64'h0 : io_vme_rd_data_bits; // @[TensorLoad.scala 236:25:@3062.4]
  assign _T_4947 = set == 4'h0; // @[TensorLoad.scala 242:51:@3093.4]
  assign _T_4948 = _T_4495 & _T_4947; // @[TensorLoad.scala 242:45:@3094.4]
  assign _T_5034 = set == 4'h1; // @[TensorLoad.scala 242:51:@3144.4]
  assign _T_5035 = _T_4495 & _T_5034; // @[TensorLoad.scala 242:45:@3145.4]
  assign _T_5121 = set == 4'h2; // @[TensorLoad.scala 242:51:@3195.4]
  assign _T_5122 = _T_4495 & _T_5121; // @[TensorLoad.scala 242:45:@3196.4]
  assign _T_5208 = set == 4'h3; // @[TensorLoad.scala 242:51:@3246.4]
  assign _T_5209 = _T_4495 & _T_5208; // @[TensorLoad.scala 242:45:@3247.4]
  assign _T_5295 = set == 4'h4; // @[TensorLoad.scala 242:51:@3297.4]
  assign _T_5296 = _T_4495 & _T_5295; // @[TensorLoad.scala 242:45:@3298.4]
  assign _T_5382 = set == 4'h5; // @[TensorLoad.scala 242:51:@3348.4]
  assign _T_5383 = _T_4495 & _T_5382; // @[TensorLoad.scala 242:45:@3349.4]
  assign _T_5469 = set == 4'h6; // @[TensorLoad.scala 242:51:@3399.4]
  assign _T_5470 = _T_4495 & _T_5469; // @[TensorLoad.scala 242:45:@3400.4]
  assign _T_5556 = set == 4'h7; // @[TensorLoad.scala 242:51:@3450.4]
  assign _T_5557 = _T_4495 & _T_5556; // @[TensorLoad.scala 242:45:@3451.4]
  assign _T_5643 = set == 4'h8; // @[TensorLoad.scala 242:51:@3501.4]
  assign _T_5644 = _T_4495 & _T_5643; // @[TensorLoad.scala 242:45:@3502.4]
  assign _T_5730 = set == 4'h9; // @[TensorLoad.scala 242:51:@3552.4]
  assign _T_5731 = _T_4495 & _T_5730; // @[TensorLoad.scala 242:45:@3553.4]
  assign _T_5817 = set == 4'ha; // @[TensorLoad.scala 242:51:@3603.4]
  assign _T_5818 = _T_4495 & _T_5817; // @[TensorLoad.scala 242:45:@3604.4]
  assign _T_5904 = set == 4'hb; // @[TensorLoad.scala 242:51:@3654.4]
  assign _T_5905 = _T_4495 & _T_5904; // @[TensorLoad.scala 242:45:@3655.4]
  assign _T_5991 = set == 4'hc; // @[TensorLoad.scala 242:51:@3705.4]
  assign _T_5992 = _T_4495 & _T_5991; // @[TensorLoad.scala 242:45:@3706.4]
  assign _T_6078 = set == 4'hd; // @[TensorLoad.scala 242:51:@3756.4]
  assign _T_6079 = _T_4495 & _T_6078; // @[TensorLoad.scala 242:45:@3757.4]
  assign _T_6165 = set == 4'he; // @[TensorLoad.scala 242:51:@3807.4]
  assign _T_6166 = _T_4495 & _T_6165; // @[TensorLoad.scala 242:45:@3808.4]
  assign _GEN_216 = io_tensor_rd_idx_valid; // @[TensorLoad.scala 256:26:@3881.4]
  assign _T_6482 = {tensorFile_0_1_rdata_0_data,tensorFile_0_0_rdata_0_data}; // @[TensorLoad.scala 259:38:@4007.4]
  assign _T_6624 = {tensorFile_1_1_rdata_1_data,tensorFile_1_0_rdata_1_data}; // @[TensorLoad.scala 259:38:@4059.4]
  assign _T_6766 = {tensorFile_2_1_rdata_2_data,tensorFile_2_0_rdata_2_data}; // @[TensorLoad.scala 259:38:@4111.4]
  assign _T_6908 = {tensorFile_3_1_rdata_3_data,tensorFile_3_0_rdata_3_data}; // @[TensorLoad.scala 259:38:@4163.4]
  assign _T_7050 = {tensorFile_4_1_rdata_4_data,tensorFile_4_0_rdata_4_data}; // @[TensorLoad.scala 259:38:@4215.4]
  assign _T_7192 = {tensorFile_5_1_rdata_5_data,tensorFile_5_0_rdata_5_data}; // @[TensorLoad.scala 259:38:@4267.4]
  assign _T_7334 = {tensorFile_6_1_rdata_6_data,tensorFile_6_0_rdata_6_data}; // @[TensorLoad.scala 259:38:@4319.4]
  assign _T_7476 = {tensorFile_7_1_rdata_7_data,tensorFile_7_0_rdata_7_data}; // @[TensorLoad.scala 259:38:@4371.4]
  assign _T_7618 = {tensorFile_8_1_rdata_8_data,tensorFile_8_0_rdata_8_data}; // @[TensorLoad.scala 259:38:@4423.4]
  assign _T_7760 = {tensorFile_9_1_rdata_9_data,tensorFile_9_0_rdata_9_data}; // @[TensorLoad.scala 259:38:@4475.4]
  assign _T_7902 = {tensorFile_10_1_rdata_10_data,tensorFile_10_0_rdata_10_data}; // @[TensorLoad.scala 259:38:@4527.4]
  assign _T_8044 = {tensorFile_11_1_rdata_11_data,tensorFile_11_0_rdata_11_data}; // @[TensorLoad.scala 259:38:@4579.4]
  assign _T_8186 = {tensorFile_12_1_rdata_12_data,tensorFile_12_0_rdata_12_data}; // @[TensorLoad.scala 259:38:@4631.4]
  assign _T_8328 = {tensorFile_13_1_rdata_13_data,tensorFile_13_0_rdata_13_data}; // @[TensorLoad.scala 259:38:@4683.4]
  assign _T_8470 = {tensorFile_14_1_rdata_14_data,tensorFile_14_0_rdata_14_data}; // @[TensorLoad.scala 259:38:@4735.4]
  assign _T_8612 = {tensorFile_15_1_rdata_15_data,tensorFile_15_0_rdata_15_data}; // @[TensorLoad.scala 259:38:@4787.4]
  assign _T_8760 = dec_ypad_1 == 4'h0; // @[TensorLoad.scala 263:96:@4843.4]
  assign done_no_pad = _T_4441 & _T_8760; // @[TensorLoad.scala 263:83:@4844.4]
  assign done_x_pad = _T_4444 & _T_8760; // @[TensorLoad.scala 264:72:@4849.4]
  assign _T_8767 = _T_4486 & dataCtrlDone; // @[TensorLoad.scala 265:37:@4851.4]
  assign done_y_pad = _T_8767 & yPadCtrl1_io_done; // @[TensorLoad.scala 265:52:@4852.4]
  assign _T_8768 = done_no_pad | done_x_pad; // @[TensorLoad.scala 266:26:@4853.4]
  assign io_done = _T_8768 | done_y_pad; // @[TensorLoad.scala 266:11:@4855.4]
  assign io_vme_rd_cmd_valid = state == 3'h3; // @[TensorLoad.scala 182:23:@2932.4]
  assign io_vme_rd_cmd_bits_addr = dataCtrl_io_addr; // @[TensorLoad.scala 183:27:@2933.4]
  assign io_vme_rd_cmd_bits_len = dataCtrl_io_len; // @[TensorLoad.scala 184:26:@2934.4]
  assign io_vme_rd_data_ready = state == 3'h4; // @[TensorLoad.scala 186:24:@2936.4]
  assign io_tensor_rd_data_valid = rvalid; // @[TensorLoad.scala 253:27:@3878.4]
  assign io_tensor_rd_data_bits_0_0 = _T_6482[7:0]; // @[TensorLoad.scala 259:33:@4043.4]
  assign io_tensor_rd_data_bits_0_1 = _T_6482[15:8]; // @[TensorLoad.scala 259:33:@4044.4]
  assign io_tensor_rd_data_bits_0_2 = _T_6482[23:16]; // @[TensorLoad.scala 259:33:@4045.4]
  assign io_tensor_rd_data_bits_0_3 = _T_6482[31:24]; // @[TensorLoad.scala 259:33:@4046.4]
  assign io_tensor_rd_data_bits_0_4 = _T_6482[39:32]; // @[TensorLoad.scala 259:33:@4047.4]
  assign io_tensor_rd_data_bits_0_5 = _T_6482[47:40]; // @[TensorLoad.scala 259:33:@4048.4]
  assign io_tensor_rd_data_bits_0_6 = _T_6482[55:48]; // @[TensorLoad.scala 259:33:@4049.4]
  assign io_tensor_rd_data_bits_0_7 = _T_6482[63:56]; // @[TensorLoad.scala 259:33:@4050.4]
  assign io_tensor_rd_data_bits_0_8 = _T_6482[71:64]; // @[TensorLoad.scala 259:33:@4051.4]
  assign io_tensor_rd_data_bits_0_9 = _T_6482[79:72]; // @[TensorLoad.scala 259:33:@4052.4]
  assign io_tensor_rd_data_bits_0_10 = _T_6482[87:80]; // @[TensorLoad.scala 259:33:@4053.4]
  assign io_tensor_rd_data_bits_0_11 = _T_6482[95:88]; // @[TensorLoad.scala 259:33:@4054.4]
  assign io_tensor_rd_data_bits_0_12 = _T_6482[103:96]; // @[TensorLoad.scala 259:33:@4055.4]
  assign io_tensor_rd_data_bits_0_13 = _T_6482[111:104]; // @[TensorLoad.scala 259:33:@4056.4]
  assign io_tensor_rd_data_bits_0_14 = _T_6482[119:112]; // @[TensorLoad.scala 259:33:@4057.4]
  assign io_tensor_rd_data_bits_0_15 = _T_6482[127:120]; // @[TensorLoad.scala 259:33:@4058.4]
  assign io_tensor_rd_data_bits_1_0 = _T_6624[7:0]; // @[TensorLoad.scala 259:33:@4095.4]
  assign io_tensor_rd_data_bits_1_1 = _T_6624[15:8]; // @[TensorLoad.scala 259:33:@4096.4]
  assign io_tensor_rd_data_bits_1_2 = _T_6624[23:16]; // @[TensorLoad.scala 259:33:@4097.4]
  assign io_tensor_rd_data_bits_1_3 = _T_6624[31:24]; // @[TensorLoad.scala 259:33:@4098.4]
  assign io_tensor_rd_data_bits_1_4 = _T_6624[39:32]; // @[TensorLoad.scala 259:33:@4099.4]
  assign io_tensor_rd_data_bits_1_5 = _T_6624[47:40]; // @[TensorLoad.scala 259:33:@4100.4]
  assign io_tensor_rd_data_bits_1_6 = _T_6624[55:48]; // @[TensorLoad.scala 259:33:@4101.4]
  assign io_tensor_rd_data_bits_1_7 = _T_6624[63:56]; // @[TensorLoad.scala 259:33:@4102.4]
  assign io_tensor_rd_data_bits_1_8 = _T_6624[71:64]; // @[TensorLoad.scala 259:33:@4103.4]
  assign io_tensor_rd_data_bits_1_9 = _T_6624[79:72]; // @[TensorLoad.scala 259:33:@4104.4]
  assign io_tensor_rd_data_bits_1_10 = _T_6624[87:80]; // @[TensorLoad.scala 259:33:@4105.4]
  assign io_tensor_rd_data_bits_1_11 = _T_6624[95:88]; // @[TensorLoad.scala 259:33:@4106.4]
  assign io_tensor_rd_data_bits_1_12 = _T_6624[103:96]; // @[TensorLoad.scala 259:33:@4107.4]
  assign io_tensor_rd_data_bits_1_13 = _T_6624[111:104]; // @[TensorLoad.scala 259:33:@4108.4]
  assign io_tensor_rd_data_bits_1_14 = _T_6624[119:112]; // @[TensorLoad.scala 259:33:@4109.4]
  assign io_tensor_rd_data_bits_1_15 = _T_6624[127:120]; // @[TensorLoad.scala 259:33:@4110.4]
  assign io_tensor_rd_data_bits_2_0 = _T_6766[7:0]; // @[TensorLoad.scala 259:33:@4147.4]
  assign io_tensor_rd_data_bits_2_1 = _T_6766[15:8]; // @[TensorLoad.scala 259:33:@4148.4]
  assign io_tensor_rd_data_bits_2_2 = _T_6766[23:16]; // @[TensorLoad.scala 259:33:@4149.4]
  assign io_tensor_rd_data_bits_2_3 = _T_6766[31:24]; // @[TensorLoad.scala 259:33:@4150.4]
  assign io_tensor_rd_data_bits_2_4 = _T_6766[39:32]; // @[TensorLoad.scala 259:33:@4151.4]
  assign io_tensor_rd_data_bits_2_5 = _T_6766[47:40]; // @[TensorLoad.scala 259:33:@4152.4]
  assign io_tensor_rd_data_bits_2_6 = _T_6766[55:48]; // @[TensorLoad.scala 259:33:@4153.4]
  assign io_tensor_rd_data_bits_2_7 = _T_6766[63:56]; // @[TensorLoad.scala 259:33:@4154.4]
  assign io_tensor_rd_data_bits_2_8 = _T_6766[71:64]; // @[TensorLoad.scala 259:33:@4155.4]
  assign io_tensor_rd_data_bits_2_9 = _T_6766[79:72]; // @[TensorLoad.scala 259:33:@4156.4]
  assign io_tensor_rd_data_bits_2_10 = _T_6766[87:80]; // @[TensorLoad.scala 259:33:@4157.4]
  assign io_tensor_rd_data_bits_2_11 = _T_6766[95:88]; // @[TensorLoad.scala 259:33:@4158.4]
  assign io_tensor_rd_data_bits_2_12 = _T_6766[103:96]; // @[TensorLoad.scala 259:33:@4159.4]
  assign io_tensor_rd_data_bits_2_13 = _T_6766[111:104]; // @[TensorLoad.scala 259:33:@4160.4]
  assign io_tensor_rd_data_bits_2_14 = _T_6766[119:112]; // @[TensorLoad.scala 259:33:@4161.4]
  assign io_tensor_rd_data_bits_2_15 = _T_6766[127:120]; // @[TensorLoad.scala 259:33:@4162.4]
  assign io_tensor_rd_data_bits_3_0 = _T_6908[7:0]; // @[TensorLoad.scala 259:33:@4199.4]
  assign io_tensor_rd_data_bits_3_1 = _T_6908[15:8]; // @[TensorLoad.scala 259:33:@4200.4]
  assign io_tensor_rd_data_bits_3_2 = _T_6908[23:16]; // @[TensorLoad.scala 259:33:@4201.4]
  assign io_tensor_rd_data_bits_3_3 = _T_6908[31:24]; // @[TensorLoad.scala 259:33:@4202.4]
  assign io_tensor_rd_data_bits_3_4 = _T_6908[39:32]; // @[TensorLoad.scala 259:33:@4203.4]
  assign io_tensor_rd_data_bits_3_5 = _T_6908[47:40]; // @[TensorLoad.scala 259:33:@4204.4]
  assign io_tensor_rd_data_bits_3_6 = _T_6908[55:48]; // @[TensorLoad.scala 259:33:@4205.4]
  assign io_tensor_rd_data_bits_3_7 = _T_6908[63:56]; // @[TensorLoad.scala 259:33:@4206.4]
  assign io_tensor_rd_data_bits_3_8 = _T_6908[71:64]; // @[TensorLoad.scala 259:33:@4207.4]
  assign io_tensor_rd_data_bits_3_9 = _T_6908[79:72]; // @[TensorLoad.scala 259:33:@4208.4]
  assign io_tensor_rd_data_bits_3_10 = _T_6908[87:80]; // @[TensorLoad.scala 259:33:@4209.4]
  assign io_tensor_rd_data_bits_3_11 = _T_6908[95:88]; // @[TensorLoad.scala 259:33:@4210.4]
  assign io_tensor_rd_data_bits_3_12 = _T_6908[103:96]; // @[TensorLoad.scala 259:33:@4211.4]
  assign io_tensor_rd_data_bits_3_13 = _T_6908[111:104]; // @[TensorLoad.scala 259:33:@4212.4]
  assign io_tensor_rd_data_bits_3_14 = _T_6908[119:112]; // @[TensorLoad.scala 259:33:@4213.4]
  assign io_tensor_rd_data_bits_3_15 = _T_6908[127:120]; // @[TensorLoad.scala 259:33:@4214.4]
  assign io_tensor_rd_data_bits_4_0 = _T_7050[7:0]; // @[TensorLoad.scala 259:33:@4251.4]
  assign io_tensor_rd_data_bits_4_1 = _T_7050[15:8]; // @[TensorLoad.scala 259:33:@4252.4]
  assign io_tensor_rd_data_bits_4_2 = _T_7050[23:16]; // @[TensorLoad.scala 259:33:@4253.4]
  assign io_tensor_rd_data_bits_4_3 = _T_7050[31:24]; // @[TensorLoad.scala 259:33:@4254.4]
  assign io_tensor_rd_data_bits_4_4 = _T_7050[39:32]; // @[TensorLoad.scala 259:33:@4255.4]
  assign io_tensor_rd_data_bits_4_5 = _T_7050[47:40]; // @[TensorLoad.scala 259:33:@4256.4]
  assign io_tensor_rd_data_bits_4_6 = _T_7050[55:48]; // @[TensorLoad.scala 259:33:@4257.4]
  assign io_tensor_rd_data_bits_4_7 = _T_7050[63:56]; // @[TensorLoad.scala 259:33:@4258.4]
  assign io_tensor_rd_data_bits_4_8 = _T_7050[71:64]; // @[TensorLoad.scala 259:33:@4259.4]
  assign io_tensor_rd_data_bits_4_9 = _T_7050[79:72]; // @[TensorLoad.scala 259:33:@4260.4]
  assign io_tensor_rd_data_bits_4_10 = _T_7050[87:80]; // @[TensorLoad.scala 259:33:@4261.4]
  assign io_tensor_rd_data_bits_4_11 = _T_7050[95:88]; // @[TensorLoad.scala 259:33:@4262.4]
  assign io_tensor_rd_data_bits_4_12 = _T_7050[103:96]; // @[TensorLoad.scala 259:33:@4263.4]
  assign io_tensor_rd_data_bits_4_13 = _T_7050[111:104]; // @[TensorLoad.scala 259:33:@4264.4]
  assign io_tensor_rd_data_bits_4_14 = _T_7050[119:112]; // @[TensorLoad.scala 259:33:@4265.4]
  assign io_tensor_rd_data_bits_4_15 = _T_7050[127:120]; // @[TensorLoad.scala 259:33:@4266.4]
  assign io_tensor_rd_data_bits_5_0 = _T_7192[7:0]; // @[TensorLoad.scala 259:33:@4303.4]
  assign io_tensor_rd_data_bits_5_1 = _T_7192[15:8]; // @[TensorLoad.scala 259:33:@4304.4]
  assign io_tensor_rd_data_bits_5_2 = _T_7192[23:16]; // @[TensorLoad.scala 259:33:@4305.4]
  assign io_tensor_rd_data_bits_5_3 = _T_7192[31:24]; // @[TensorLoad.scala 259:33:@4306.4]
  assign io_tensor_rd_data_bits_5_4 = _T_7192[39:32]; // @[TensorLoad.scala 259:33:@4307.4]
  assign io_tensor_rd_data_bits_5_5 = _T_7192[47:40]; // @[TensorLoad.scala 259:33:@4308.4]
  assign io_tensor_rd_data_bits_5_6 = _T_7192[55:48]; // @[TensorLoad.scala 259:33:@4309.4]
  assign io_tensor_rd_data_bits_5_7 = _T_7192[63:56]; // @[TensorLoad.scala 259:33:@4310.4]
  assign io_tensor_rd_data_bits_5_8 = _T_7192[71:64]; // @[TensorLoad.scala 259:33:@4311.4]
  assign io_tensor_rd_data_bits_5_9 = _T_7192[79:72]; // @[TensorLoad.scala 259:33:@4312.4]
  assign io_tensor_rd_data_bits_5_10 = _T_7192[87:80]; // @[TensorLoad.scala 259:33:@4313.4]
  assign io_tensor_rd_data_bits_5_11 = _T_7192[95:88]; // @[TensorLoad.scala 259:33:@4314.4]
  assign io_tensor_rd_data_bits_5_12 = _T_7192[103:96]; // @[TensorLoad.scala 259:33:@4315.4]
  assign io_tensor_rd_data_bits_5_13 = _T_7192[111:104]; // @[TensorLoad.scala 259:33:@4316.4]
  assign io_tensor_rd_data_bits_5_14 = _T_7192[119:112]; // @[TensorLoad.scala 259:33:@4317.4]
  assign io_tensor_rd_data_bits_5_15 = _T_7192[127:120]; // @[TensorLoad.scala 259:33:@4318.4]
  assign io_tensor_rd_data_bits_6_0 = _T_7334[7:0]; // @[TensorLoad.scala 259:33:@4355.4]
  assign io_tensor_rd_data_bits_6_1 = _T_7334[15:8]; // @[TensorLoad.scala 259:33:@4356.4]
  assign io_tensor_rd_data_bits_6_2 = _T_7334[23:16]; // @[TensorLoad.scala 259:33:@4357.4]
  assign io_tensor_rd_data_bits_6_3 = _T_7334[31:24]; // @[TensorLoad.scala 259:33:@4358.4]
  assign io_tensor_rd_data_bits_6_4 = _T_7334[39:32]; // @[TensorLoad.scala 259:33:@4359.4]
  assign io_tensor_rd_data_bits_6_5 = _T_7334[47:40]; // @[TensorLoad.scala 259:33:@4360.4]
  assign io_tensor_rd_data_bits_6_6 = _T_7334[55:48]; // @[TensorLoad.scala 259:33:@4361.4]
  assign io_tensor_rd_data_bits_6_7 = _T_7334[63:56]; // @[TensorLoad.scala 259:33:@4362.4]
  assign io_tensor_rd_data_bits_6_8 = _T_7334[71:64]; // @[TensorLoad.scala 259:33:@4363.4]
  assign io_tensor_rd_data_bits_6_9 = _T_7334[79:72]; // @[TensorLoad.scala 259:33:@4364.4]
  assign io_tensor_rd_data_bits_6_10 = _T_7334[87:80]; // @[TensorLoad.scala 259:33:@4365.4]
  assign io_tensor_rd_data_bits_6_11 = _T_7334[95:88]; // @[TensorLoad.scala 259:33:@4366.4]
  assign io_tensor_rd_data_bits_6_12 = _T_7334[103:96]; // @[TensorLoad.scala 259:33:@4367.4]
  assign io_tensor_rd_data_bits_6_13 = _T_7334[111:104]; // @[TensorLoad.scala 259:33:@4368.4]
  assign io_tensor_rd_data_bits_6_14 = _T_7334[119:112]; // @[TensorLoad.scala 259:33:@4369.4]
  assign io_tensor_rd_data_bits_6_15 = _T_7334[127:120]; // @[TensorLoad.scala 259:33:@4370.4]
  assign io_tensor_rd_data_bits_7_0 = _T_7476[7:0]; // @[TensorLoad.scala 259:33:@4407.4]
  assign io_tensor_rd_data_bits_7_1 = _T_7476[15:8]; // @[TensorLoad.scala 259:33:@4408.4]
  assign io_tensor_rd_data_bits_7_2 = _T_7476[23:16]; // @[TensorLoad.scala 259:33:@4409.4]
  assign io_tensor_rd_data_bits_7_3 = _T_7476[31:24]; // @[TensorLoad.scala 259:33:@4410.4]
  assign io_tensor_rd_data_bits_7_4 = _T_7476[39:32]; // @[TensorLoad.scala 259:33:@4411.4]
  assign io_tensor_rd_data_bits_7_5 = _T_7476[47:40]; // @[TensorLoad.scala 259:33:@4412.4]
  assign io_tensor_rd_data_bits_7_6 = _T_7476[55:48]; // @[TensorLoad.scala 259:33:@4413.4]
  assign io_tensor_rd_data_bits_7_7 = _T_7476[63:56]; // @[TensorLoad.scala 259:33:@4414.4]
  assign io_tensor_rd_data_bits_7_8 = _T_7476[71:64]; // @[TensorLoad.scala 259:33:@4415.4]
  assign io_tensor_rd_data_bits_7_9 = _T_7476[79:72]; // @[TensorLoad.scala 259:33:@4416.4]
  assign io_tensor_rd_data_bits_7_10 = _T_7476[87:80]; // @[TensorLoad.scala 259:33:@4417.4]
  assign io_tensor_rd_data_bits_7_11 = _T_7476[95:88]; // @[TensorLoad.scala 259:33:@4418.4]
  assign io_tensor_rd_data_bits_7_12 = _T_7476[103:96]; // @[TensorLoad.scala 259:33:@4419.4]
  assign io_tensor_rd_data_bits_7_13 = _T_7476[111:104]; // @[TensorLoad.scala 259:33:@4420.4]
  assign io_tensor_rd_data_bits_7_14 = _T_7476[119:112]; // @[TensorLoad.scala 259:33:@4421.4]
  assign io_tensor_rd_data_bits_7_15 = _T_7476[127:120]; // @[TensorLoad.scala 259:33:@4422.4]
  assign io_tensor_rd_data_bits_8_0 = _T_7618[7:0]; // @[TensorLoad.scala 259:33:@4459.4]
  assign io_tensor_rd_data_bits_8_1 = _T_7618[15:8]; // @[TensorLoad.scala 259:33:@4460.4]
  assign io_tensor_rd_data_bits_8_2 = _T_7618[23:16]; // @[TensorLoad.scala 259:33:@4461.4]
  assign io_tensor_rd_data_bits_8_3 = _T_7618[31:24]; // @[TensorLoad.scala 259:33:@4462.4]
  assign io_tensor_rd_data_bits_8_4 = _T_7618[39:32]; // @[TensorLoad.scala 259:33:@4463.4]
  assign io_tensor_rd_data_bits_8_5 = _T_7618[47:40]; // @[TensorLoad.scala 259:33:@4464.4]
  assign io_tensor_rd_data_bits_8_6 = _T_7618[55:48]; // @[TensorLoad.scala 259:33:@4465.4]
  assign io_tensor_rd_data_bits_8_7 = _T_7618[63:56]; // @[TensorLoad.scala 259:33:@4466.4]
  assign io_tensor_rd_data_bits_8_8 = _T_7618[71:64]; // @[TensorLoad.scala 259:33:@4467.4]
  assign io_tensor_rd_data_bits_8_9 = _T_7618[79:72]; // @[TensorLoad.scala 259:33:@4468.4]
  assign io_tensor_rd_data_bits_8_10 = _T_7618[87:80]; // @[TensorLoad.scala 259:33:@4469.4]
  assign io_tensor_rd_data_bits_8_11 = _T_7618[95:88]; // @[TensorLoad.scala 259:33:@4470.4]
  assign io_tensor_rd_data_bits_8_12 = _T_7618[103:96]; // @[TensorLoad.scala 259:33:@4471.4]
  assign io_tensor_rd_data_bits_8_13 = _T_7618[111:104]; // @[TensorLoad.scala 259:33:@4472.4]
  assign io_tensor_rd_data_bits_8_14 = _T_7618[119:112]; // @[TensorLoad.scala 259:33:@4473.4]
  assign io_tensor_rd_data_bits_8_15 = _T_7618[127:120]; // @[TensorLoad.scala 259:33:@4474.4]
  assign io_tensor_rd_data_bits_9_0 = _T_7760[7:0]; // @[TensorLoad.scala 259:33:@4511.4]
  assign io_tensor_rd_data_bits_9_1 = _T_7760[15:8]; // @[TensorLoad.scala 259:33:@4512.4]
  assign io_tensor_rd_data_bits_9_2 = _T_7760[23:16]; // @[TensorLoad.scala 259:33:@4513.4]
  assign io_tensor_rd_data_bits_9_3 = _T_7760[31:24]; // @[TensorLoad.scala 259:33:@4514.4]
  assign io_tensor_rd_data_bits_9_4 = _T_7760[39:32]; // @[TensorLoad.scala 259:33:@4515.4]
  assign io_tensor_rd_data_bits_9_5 = _T_7760[47:40]; // @[TensorLoad.scala 259:33:@4516.4]
  assign io_tensor_rd_data_bits_9_6 = _T_7760[55:48]; // @[TensorLoad.scala 259:33:@4517.4]
  assign io_tensor_rd_data_bits_9_7 = _T_7760[63:56]; // @[TensorLoad.scala 259:33:@4518.4]
  assign io_tensor_rd_data_bits_9_8 = _T_7760[71:64]; // @[TensorLoad.scala 259:33:@4519.4]
  assign io_tensor_rd_data_bits_9_9 = _T_7760[79:72]; // @[TensorLoad.scala 259:33:@4520.4]
  assign io_tensor_rd_data_bits_9_10 = _T_7760[87:80]; // @[TensorLoad.scala 259:33:@4521.4]
  assign io_tensor_rd_data_bits_9_11 = _T_7760[95:88]; // @[TensorLoad.scala 259:33:@4522.4]
  assign io_tensor_rd_data_bits_9_12 = _T_7760[103:96]; // @[TensorLoad.scala 259:33:@4523.4]
  assign io_tensor_rd_data_bits_9_13 = _T_7760[111:104]; // @[TensorLoad.scala 259:33:@4524.4]
  assign io_tensor_rd_data_bits_9_14 = _T_7760[119:112]; // @[TensorLoad.scala 259:33:@4525.4]
  assign io_tensor_rd_data_bits_9_15 = _T_7760[127:120]; // @[TensorLoad.scala 259:33:@4526.4]
  assign io_tensor_rd_data_bits_10_0 = _T_7902[7:0]; // @[TensorLoad.scala 259:33:@4563.4]
  assign io_tensor_rd_data_bits_10_1 = _T_7902[15:8]; // @[TensorLoad.scala 259:33:@4564.4]
  assign io_tensor_rd_data_bits_10_2 = _T_7902[23:16]; // @[TensorLoad.scala 259:33:@4565.4]
  assign io_tensor_rd_data_bits_10_3 = _T_7902[31:24]; // @[TensorLoad.scala 259:33:@4566.4]
  assign io_tensor_rd_data_bits_10_4 = _T_7902[39:32]; // @[TensorLoad.scala 259:33:@4567.4]
  assign io_tensor_rd_data_bits_10_5 = _T_7902[47:40]; // @[TensorLoad.scala 259:33:@4568.4]
  assign io_tensor_rd_data_bits_10_6 = _T_7902[55:48]; // @[TensorLoad.scala 259:33:@4569.4]
  assign io_tensor_rd_data_bits_10_7 = _T_7902[63:56]; // @[TensorLoad.scala 259:33:@4570.4]
  assign io_tensor_rd_data_bits_10_8 = _T_7902[71:64]; // @[TensorLoad.scala 259:33:@4571.4]
  assign io_tensor_rd_data_bits_10_9 = _T_7902[79:72]; // @[TensorLoad.scala 259:33:@4572.4]
  assign io_tensor_rd_data_bits_10_10 = _T_7902[87:80]; // @[TensorLoad.scala 259:33:@4573.4]
  assign io_tensor_rd_data_bits_10_11 = _T_7902[95:88]; // @[TensorLoad.scala 259:33:@4574.4]
  assign io_tensor_rd_data_bits_10_12 = _T_7902[103:96]; // @[TensorLoad.scala 259:33:@4575.4]
  assign io_tensor_rd_data_bits_10_13 = _T_7902[111:104]; // @[TensorLoad.scala 259:33:@4576.4]
  assign io_tensor_rd_data_bits_10_14 = _T_7902[119:112]; // @[TensorLoad.scala 259:33:@4577.4]
  assign io_tensor_rd_data_bits_10_15 = _T_7902[127:120]; // @[TensorLoad.scala 259:33:@4578.4]
  assign io_tensor_rd_data_bits_11_0 = _T_8044[7:0]; // @[TensorLoad.scala 259:33:@4615.4]
  assign io_tensor_rd_data_bits_11_1 = _T_8044[15:8]; // @[TensorLoad.scala 259:33:@4616.4]
  assign io_tensor_rd_data_bits_11_2 = _T_8044[23:16]; // @[TensorLoad.scala 259:33:@4617.4]
  assign io_tensor_rd_data_bits_11_3 = _T_8044[31:24]; // @[TensorLoad.scala 259:33:@4618.4]
  assign io_tensor_rd_data_bits_11_4 = _T_8044[39:32]; // @[TensorLoad.scala 259:33:@4619.4]
  assign io_tensor_rd_data_bits_11_5 = _T_8044[47:40]; // @[TensorLoad.scala 259:33:@4620.4]
  assign io_tensor_rd_data_bits_11_6 = _T_8044[55:48]; // @[TensorLoad.scala 259:33:@4621.4]
  assign io_tensor_rd_data_bits_11_7 = _T_8044[63:56]; // @[TensorLoad.scala 259:33:@4622.4]
  assign io_tensor_rd_data_bits_11_8 = _T_8044[71:64]; // @[TensorLoad.scala 259:33:@4623.4]
  assign io_tensor_rd_data_bits_11_9 = _T_8044[79:72]; // @[TensorLoad.scala 259:33:@4624.4]
  assign io_tensor_rd_data_bits_11_10 = _T_8044[87:80]; // @[TensorLoad.scala 259:33:@4625.4]
  assign io_tensor_rd_data_bits_11_11 = _T_8044[95:88]; // @[TensorLoad.scala 259:33:@4626.4]
  assign io_tensor_rd_data_bits_11_12 = _T_8044[103:96]; // @[TensorLoad.scala 259:33:@4627.4]
  assign io_tensor_rd_data_bits_11_13 = _T_8044[111:104]; // @[TensorLoad.scala 259:33:@4628.4]
  assign io_tensor_rd_data_bits_11_14 = _T_8044[119:112]; // @[TensorLoad.scala 259:33:@4629.4]
  assign io_tensor_rd_data_bits_11_15 = _T_8044[127:120]; // @[TensorLoad.scala 259:33:@4630.4]
  assign io_tensor_rd_data_bits_12_0 = _T_8186[7:0]; // @[TensorLoad.scala 259:33:@4667.4]
  assign io_tensor_rd_data_bits_12_1 = _T_8186[15:8]; // @[TensorLoad.scala 259:33:@4668.4]
  assign io_tensor_rd_data_bits_12_2 = _T_8186[23:16]; // @[TensorLoad.scala 259:33:@4669.4]
  assign io_tensor_rd_data_bits_12_3 = _T_8186[31:24]; // @[TensorLoad.scala 259:33:@4670.4]
  assign io_tensor_rd_data_bits_12_4 = _T_8186[39:32]; // @[TensorLoad.scala 259:33:@4671.4]
  assign io_tensor_rd_data_bits_12_5 = _T_8186[47:40]; // @[TensorLoad.scala 259:33:@4672.4]
  assign io_tensor_rd_data_bits_12_6 = _T_8186[55:48]; // @[TensorLoad.scala 259:33:@4673.4]
  assign io_tensor_rd_data_bits_12_7 = _T_8186[63:56]; // @[TensorLoad.scala 259:33:@4674.4]
  assign io_tensor_rd_data_bits_12_8 = _T_8186[71:64]; // @[TensorLoad.scala 259:33:@4675.4]
  assign io_tensor_rd_data_bits_12_9 = _T_8186[79:72]; // @[TensorLoad.scala 259:33:@4676.4]
  assign io_tensor_rd_data_bits_12_10 = _T_8186[87:80]; // @[TensorLoad.scala 259:33:@4677.4]
  assign io_tensor_rd_data_bits_12_11 = _T_8186[95:88]; // @[TensorLoad.scala 259:33:@4678.4]
  assign io_tensor_rd_data_bits_12_12 = _T_8186[103:96]; // @[TensorLoad.scala 259:33:@4679.4]
  assign io_tensor_rd_data_bits_12_13 = _T_8186[111:104]; // @[TensorLoad.scala 259:33:@4680.4]
  assign io_tensor_rd_data_bits_12_14 = _T_8186[119:112]; // @[TensorLoad.scala 259:33:@4681.4]
  assign io_tensor_rd_data_bits_12_15 = _T_8186[127:120]; // @[TensorLoad.scala 259:33:@4682.4]
  assign io_tensor_rd_data_bits_13_0 = _T_8328[7:0]; // @[TensorLoad.scala 259:33:@4719.4]
  assign io_tensor_rd_data_bits_13_1 = _T_8328[15:8]; // @[TensorLoad.scala 259:33:@4720.4]
  assign io_tensor_rd_data_bits_13_2 = _T_8328[23:16]; // @[TensorLoad.scala 259:33:@4721.4]
  assign io_tensor_rd_data_bits_13_3 = _T_8328[31:24]; // @[TensorLoad.scala 259:33:@4722.4]
  assign io_tensor_rd_data_bits_13_4 = _T_8328[39:32]; // @[TensorLoad.scala 259:33:@4723.4]
  assign io_tensor_rd_data_bits_13_5 = _T_8328[47:40]; // @[TensorLoad.scala 259:33:@4724.4]
  assign io_tensor_rd_data_bits_13_6 = _T_8328[55:48]; // @[TensorLoad.scala 259:33:@4725.4]
  assign io_tensor_rd_data_bits_13_7 = _T_8328[63:56]; // @[TensorLoad.scala 259:33:@4726.4]
  assign io_tensor_rd_data_bits_13_8 = _T_8328[71:64]; // @[TensorLoad.scala 259:33:@4727.4]
  assign io_tensor_rd_data_bits_13_9 = _T_8328[79:72]; // @[TensorLoad.scala 259:33:@4728.4]
  assign io_tensor_rd_data_bits_13_10 = _T_8328[87:80]; // @[TensorLoad.scala 259:33:@4729.4]
  assign io_tensor_rd_data_bits_13_11 = _T_8328[95:88]; // @[TensorLoad.scala 259:33:@4730.4]
  assign io_tensor_rd_data_bits_13_12 = _T_8328[103:96]; // @[TensorLoad.scala 259:33:@4731.4]
  assign io_tensor_rd_data_bits_13_13 = _T_8328[111:104]; // @[TensorLoad.scala 259:33:@4732.4]
  assign io_tensor_rd_data_bits_13_14 = _T_8328[119:112]; // @[TensorLoad.scala 259:33:@4733.4]
  assign io_tensor_rd_data_bits_13_15 = _T_8328[127:120]; // @[TensorLoad.scala 259:33:@4734.4]
  assign io_tensor_rd_data_bits_14_0 = _T_8470[7:0]; // @[TensorLoad.scala 259:33:@4771.4]
  assign io_tensor_rd_data_bits_14_1 = _T_8470[15:8]; // @[TensorLoad.scala 259:33:@4772.4]
  assign io_tensor_rd_data_bits_14_2 = _T_8470[23:16]; // @[TensorLoad.scala 259:33:@4773.4]
  assign io_tensor_rd_data_bits_14_3 = _T_8470[31:24]; // @[TensorLoad.scala 259:33:@4774.4]
  assign io_tensor_rd_data_bits_14_4 = _T_8470[39:32]; // @[TensorLoad.scala 259:33:@4775.4]
  assign io_tensor_rd_data_bits_14_5 = _T_8470[47:40]; // @[TensorLoad.scala 259:33:@4776.4]
  assign io_tensor_rd_data_bits_14_6 = _T_8470[55:48]; // @[TensorLoad.scala 259:33:@4777.4]
  assign io_tensor_rd_data_bits_14_7 = _T_8470[63:56]; // @[TensorLoad.scala 259:33:@4778.4]
  assign io_tensor_rd_data_bits_14_8 = _T_8470[71:64]; // @[TensorLoad.scala 259:33:@4779.4]
  assign io_tensor_rd_data_bits_14_9 = _T_8470[79:72]; // @[TensorLoad.scala 259:33:@4780.4]
  assign io_tensor_rd_data_bits_14_10 = _T_8470[87:80]; // @[TensorLoad.scala 259:33:@4781.4]
  assign io_tensor_rd_data_bits_14_11 = _T_8470[95:88]; // @[TensorLoad.scala 259:33:@4782.4]
  assign io_tensor_rd_data_bits_14_12 = _T_8470[103:96]; // @[TensorLoad.scala 259:33:@4783.4]
  assign io_tensor_rd_data_bits_14_13 = _T_8470[111:104]; // @[TensorLoad.scala 259:33:@4784.4]
  assign io_tensor_rd_data_bits_14_14 = _T_8470[119:112]; // @[TensorLoad.scala 259:33:@4785.4]
  assign io_tensor_rd_data_bits_14_15 = _T_8470[127:120]; // @[TensorLoad.scala 259:33:@4786.4]
  assign io_tensor_rd_data_bits_15_0 = _T_8612[7:0]; // @[TensorLoad.scala 259:33:@4823.4]
  assign io_tensor_rd_data_bits_15_1 = _T_8612[15:8]; // @[TensorLoad.scala 259:33:@4824.4]
  assign io_tensor_rd_data_bits_15_2 = _T_8612[23:16]; // @[TensorLoad.scala 259:33:@4825.4]
  assign io_tensor_rd_data_bits_15_3 = _T_8612[31:24]; // @[TensorLoad.scala 259:33:@4826.4]
  assign io_tensor_rd_data_bits_15_4 = _T_8612[39:32]; // @[TensorLoad.scala 259:33:@4827.4]
  assign io_tensor_rd_data_bits_15_5 = _T_8612[47:40]; // @[TensorLoad.scala 259:33:@4828.4]
  assign io_tensor_rd_data_bits_15_6 = _T_8612[55:48]; // @[TensorLoad.scala 259:33:@4829.4]
  assign io_tensor_rd_data_bits_15_7 = _T_8612[63:56]; // @[TensorLoad.scala 259:33:@4830.4]
  assign io_tensor_rd_data_bits_15_8 = _T_8612[71:64]; // @[TensorLoad.scala 259:33:@4831.4]
  assign io_tensor_rd_data_bits_15_9 = _T_8612[79:72]; // @[TensorLoad.scala 259:33:@4832.4]
  assign io_tensor_rd_data_bits_15_10 = _T_8612[87:80]; // @[TensorLoad.scala 259:33:@4833.4]
  assign io_tensor_rd_data_bits_15_11 = _T_8612[95:88]; // @[TensorLoad.scala 259:33:@4834.4]
  assign io_tensor_rd_data_bits_15_12 = _T_8612[103:96]; // @[TensorLoad.scala 259:33:@4835.4]
  assign io_tensor_rd_data_bits_15_13 = _T_8612[111:104]; // @[TensorLoad.scala 259:33:@4836.4]
  assign io_tensor_rd_data_bits_15_14 = _T_8612[119:112]; // @[TensorLoad.scala 259:33:@4837.4]
  assign io_tensor_rd_data_bits_15_15 = _T_8612[127:120]; // @[TensorLoad.scala 259:33:@4838.4]
  assign dataCtrl_clock = clock; // @[:@2727.4]
  assign dataCtrl_io_start = _T_4420 & io_start; // @[TensorLoad.scala 147:21:@2862.4]
  assign dataCtrl_io_inst = io_inst; // @[TensorLoad.scala 148:20:@2863.4]
  assign dataCtrl_io_baddr = io_baddr; // @[TensorLoad.scala 149:21:@2864.4]
  assign dataCtrl_io_xinit = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[TensorLoad.scala 150:21:@2866.4]
  assign dataCtrl_io_xupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 151:23:@2868.4]
  assign dataCtrl_io_yupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 152:23:@2870.4]
  assign yPadCtrl0_clock = clock; // @[:@2731.4]
  assign yPadCtrl0_reset = reset; // @[:@2732.4]
  assign yPadCtrl0_io_start = _T_4433 & io_start; // @[TensorLoad.scala 161:22:@2885.4]
  assign yPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 176:21:@2927.4]
  assign yPadCtrl1_clock = clock; // @[:@2734.4]
  assign yPadCtrl1_reset = reset; // @[:@2735.4]
  assign yPadCtrl1_io_start = _T_4408 & _T_4445; // @[TensorLoad.scala 163:22:@2896.4]
  assign yPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 177:21:@2928.4]
  assign xPadCtrl0_clock = clock; // @[:@2737.4]
  assign xPadCtrl0_reset = reset; // @[:@2738.4]
  assign xPadCtrl0_io_start = _T_4398 & _T_4466; // @[TensorLoad.scala 167:22:@2916.4]
  assign xPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 178:21:@2929.4]
  assign xPadCtrl1_clock = clock; // @[:@2740.4]
  assign xPadCtrl1_reset = reset; // @[:@2741.4]
  assign xPadCtrl1_io_start = _T_4471 & _T_4477; // @[TensorLoad.scala 173:22:@2926.4]
  assign xPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 179:21:@2930.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_0_0[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_0_1[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_1_0[initvar] = _RAND_2[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_1_1[initvar] = _RAND_3[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_2_0[initvar] = _RAND_4[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_2_1[initvar] = _RAND_5[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_3_0[initvar] = _RAND_6[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_3_1[initvar] = _RAND_7[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_4_0[initvar] = _RAND_8[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_4_1[initvar] = _RAND_9[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_5_0[initvar] = _RAND_10[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_5_1[initvar] = _RAND_11[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_12 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_6_0[initvar] = _RAND_12[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_6_1[initvar] = _RAND_13[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_14 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_7_0[initvar] = _RAND_14[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_15 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_7_1[initvar] = _RAND_15[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_16 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_8_0[initvar] = _RAND_16[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_8_1[initvar] = _RAND_17[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_18 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_9_0[initvar] = _RAND_18[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_19 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_9_1[initvar] = _RAND_19[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_20 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_10_0[initvar] = _RAND_20[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_10_1[initvar] = _RAND_21[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_22 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_11_0[initvar] = _RAND_22[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_23 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_11_1[initvar] = _RAND_23[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_24 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_12_0[initvar] = _RAND_24[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_12_1[initvar] = _RAND_25[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_26 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_13_0[initvar] = _RAND_26[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_27 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_13_1[initvar] = _RAND_27[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_28 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_14_0[initvar] = _RAND_28[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_14_1[initvar] = _RAND_29[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_30 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_15_0[initvar] = _RAND_30[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_31 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_15_1[initvar] = _RAND_31[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  dataCtrlDone = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  tag = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  set = _RAND_34[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  state = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  waddr_cur = _RAND_36[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  waddr_nxt = _RAND_37[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  rvalid = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  tensorFile_0_0_rdata_0_addr_pipe_0 = _RAND_39[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  tensorFile_0_1_rdata_0_addr_pipe_0 = _RAND_40[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  tensorFile_1_0_rdata_1_addr_pipe_0 = _RAND_41[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  tensorFile_1_1_rdata_1_addr_pipe_0 = _RAND_42[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  tensorFile_2_0_rdata_2_addr_pipe_0 = _RAND_43[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  tensorFile_2_1_rdata_2_addr_pipe_0 = _RAND_44[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  tensorFile_3_0_rdata_3_addr_pipe_0 = _RAND_45[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  tensorFile_3_1_rdata_3_addr_pipe_0 = _RAND_46[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  tensorFile_4_0_rdata_4_addr_pipe_0 = _RAND_47[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  tensorFile_4_1_rdata_4_addr_pipe_0 = _RAND_48[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  tensorFile_5_0_rdata_5_addr_pipe_0 = _RAND_49[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  tensorFile_5_1_rdata_5_addr_pipe_0 = _RAND_50[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  tensorFile_6_0_rdata_6_addr_pipe_0 = _RAND_51[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  tensorFile_6_1_rdata_6_addr_pipe_0 = _RAND_52[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  tensorFile_7_0_rdata_7_addr_pipe_0 = _RAND_53[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  tensorFile_7_1_rdata_7_addr_pipe_0 = _RAND_54[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  tensorFile_8_0_rdata_8_addr_pipe_0 = _RAND_55[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  tensorFile_8_1_rdata_8_addr_pipe_0 = _RAND_56[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  tensorFile_9_0_rdata_9_addr_pipe_0 = _RAND_57[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  tensorFile_9_1_rdata_9_addr_pipe_0 = _RAND_58[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  tensorFile_10_0_rdata_10_addr_pipe_0 = _RAND_59[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  tensorFile_10_1_rdata_10_addr_pipe_0 = _RAND_60[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  tensorFile_11_0_rdata_11_addr_pipe_0 = _RAND_61[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  tensorFile_11_1_rdata_11_addr_pipe_0 = _RAND_62[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  tensorFile_12_0_rdata_12_addr_pipe_0 = _RAND_63[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  tensorFile_12_1_rdata_12_addr_pipe_0 = _RAND_64[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  tensorFile_13_0_rdata_13_addr_pipe_0 = _RAND_65[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  tensorFile_13_1_rdata_13_addr_pipe_0 = _RAND_66[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  tensorFile_14_0_rdata_14_addr_pipe_0 = _RAND_67[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  tensorFile_14_1_rdata_14_addr_pipe_0 = _RAND_68[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  tensorFile_15_0_rdata_15_addr_pipe_0 = _RAND_69[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  tensorFile_15_1_rdata_15_addr_pipe_0 = _RAND_70[9:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tensorFile_0_0__T_4976_en & tensorFile_0_0__T_4976_mask) begin
      tensorFile_0_0[tensorFile_0_0__T_4976_addr] <= tensorFile_0_0__T_4976_data; // @[TensorLoad.scala 222:16:@3009.4]
    end
    if(tensorFile_0_1__T_4976_en & tensorFile_0_1__T_4976_mask) begin
      tensorFile_0_1[tensorFile_0_1__T_4976_addr] <= tensorFile_0_1__T_4976_data; // @[TensorLoad.scala 222:16:@3009.4]
    end
    if(tensorFile_1_0__T_5063_en & tensorFile_1_0__T_5063_mask) begin
      tensorFile_1_0[tensorFile_1_0__T_5063_addr] <= tensorFile_1_0__T_5063_data; // @[TensorLoad.scala 222:16:@3010.4]
    end
    if(tensorFile_1_1__T_5063_en & tensorFile_1_1__T_5063_mask) begin
      tensorFile_1_1[tensorFile_1_1__T_5063_addr] <= tensorFile_1_1__T_5063_data; // @[TensorLoad.scala 222:16:@3010.4]
    end
    if(tensorFile_2_0__T_5150_en & tensorFile_2_0__T_5150_mask) begin
      tensorFile_2_0[tensorFile_2_0__T_5150_addr] <= tensorFile_2_0__T_5150_data; // @[TensorLoad.scala 222:16:@3011.4]
    end
    if(tensorFile_2_1__T_5150_en & tensorFile_2_1__T_5150_mask) begin
      tensorFile_2_1[tensorFile_2_1__T_5150_addr] <= tensorFile_2_1__T_5150_data; // @[TensorLoad.scala 222:16:@3011.4]
    end
    if(tensorFile_3_0__T_5237_en & tensorFile_3_0__T_5237_mask) begin
      tensorFile_3_0[tensorFile_3_0__T_5237_addr] <= tensorFile_3_0__T_5237_data; // @[TensorLoad.scala 222:16:@3012.4]
    end
    if(tensorFile_3_1__T_5237_en & tensorFile_3_1__T_5237_mask) begin
      tensorFile_3_1[tensorFile_3_1__T_5237_addr] <= tensorFile_3_1__T_5237_data; // @[TensorLoad.scala 222:16:@3012.4]
    end
    if(tensorFile_4_0__T_5324_en & tensorFile_4_0__T_5324_mask) begin
      tensorFile_4_0[tensorFile_4_0__T_5324_addr] <= tensorFile_4_0__T_5324_data; // @[TensorLoad.scala 222:16:@3013.4]
    end
    if(tensorFile_4_1__T_5324_en & tensorFile_4_1__T_5324_mask) begin
      tensorFile_4_1[tensorFile_4_1__T_5324_addr] <= tensorFile_4_1__T_5324_data; // @[TensorLoad.scala 222:16:@3013.4]
    end
    if(tensorFile_5_0__T_5411_en & tensorFile_5_0__T_5411_mask) begin
      tensorFile_5_0[tensorFile_5_0__T_5411_addr] <= tensorFile_5_0__T_5411_data; // @[TensorLoad.scala 222:16:@3014.4]
    end
    if(tensorFile_5_1__T_5411_en & tensorFile_5_1__T_5411_mask) begin
      tensorFile_5_1[tensorFile_5_1__T_5411_addr] <= tensorFile_5_1__T_5411_data; // @[TensorLoad.scala 222:16:@3014.4]
    end
    if(tensorFile_6_0__T_5498_en & tensorFile_6_0__T_5498_mask) begin
      tensorFile_6_0[tensorFile_6_0__T_5498_addr] <= tensorFile_6_0__T_5498_data; // @[TensorLoad.scala 222:16:@3015.4]
    end
    if(tensorFile_6_1__T_5498_en & tensorFile_6_1__T_5498_mask) begin
      tensorFile_6_1[tensorFile_6_1__T_5498_addr] <= tensorFile_6_1__T_5498_data; // @[TensorLoad.scala 222:16:@3015.4]
    end
    if(tensorFile_7_0__T_5585_en & tensorFile_7_0__T_5585_mask) begin
      tensorFile_7_0[tensorFile_7_0__T_5585_addr] <= tensorFile_7_0__T_5585_data; // @[TensorLoad.scala 222:16:@3016.4]
    end
    if(tensorFile_7_1__T_5585_en & tensorFile_7_1__T_5585_mask) begin
      tensorFile_7_1[tensorFile_7_1__T_5585_addr] <= tensorFile_7_1__T_5585_data; // @[TensorLoad.scala 222:16:@3016.4]
    end
    if(tensorFile_8_0__T_5672_en & tensorFile_8_0__T_5672_mask) begin
      tensorFile_8_0[tensorFile_8_0__T_5672_addr] <= tensorFile_8_0__T_5672_data; // @[TensorLoad.scala 222:16:@3017.4]
    end
    if(tensorFile_8_1__T_5672_en & tensorFile_8_1__T_5672_mask) begin
      tensorFile_8_1[tensorFile_8_1__T_5672_addr] <= tensorFile_8_1__T_5672_data; // @[TensorLoad.scala 222:16:@3017.4]
    end
    if(tensorFile_9_0__T_5759_en & tensorFile_9_0__T_5759_mask) begin
      tensorFile_9_0[tensorFile_9_0__T_5759_addr] <= tensorFile_9_0__T_5759_data; // @[TensorLoad.scala 222:16:@3018.4]
    end
    if(tensorFile_9_1__T_5759_en & tensorFile_9_1__T_5759_mask) begin
      tensorFile_9_1[tensorFile_9_1__T_5759_addr] <= tensorFile_9_1__T_5759_data; // @[TensorLoad.scala 222:16:@3018.4]
    end
    if(tensorFile_10_0__T_5846_en & tensorFile_10_0__T_5846_mask) begin
      tensorFile_10_0[tensorFile_10_0__T_5846_addr] <= tensorFile_10_0__T_5846_data; // @[TensorLoad.scala 222:16:@3019.4]
    end
    if(tensorFile_10_1__T_5846_en & tensorFile_10_1__T_5846_mask) begin
      tensorFile_10_1[tensorFile_10_1__T_5846_addr] <= tensorFile_10_1__T_5846_data; // @[TensorLoad.scala 222:16:@3019.4]
    end
    if(tensorFile_11_0__T_5933_en & tensorFile_11_0__T_5933_mask) begin
      tensorFile_11_0[tensorFile_11_0__T_5933_addr] <= tensorFile_11_0__T_5933_data; // @[TensorLoad.scala 222:16:@3020.4]
    end
    if(tensorFile_11_1__T_5933_en & tensorFile_11_1__T_5933_mask) begin
      tensorFile_11_1[tensorFile_11_1__T_5933_addr] <= tensorFile_11_1__T_5933_data; // @[TensorLoad.scala 222:16:@3020.4]
    end
    if(tensorFile_12_0__T_6020_en & tensorFile_12_0__T_6020_mask) begin
      tensorFile_12_0[tensorFile_12_0__T_6020_addr] <= tensorFile_12_0__T_6020_data; // @[TensorLoad.scala 222:16:@3021.4]
    end
    if(tensorFile_12_1__T_6020_en & tensorFile_12_1__T_6020_mask) begin
      tensorFile_12_1[tensorFile_12_1__T_6020_addr] <= tensorFile_12_1__T_6020_data; // @[TensorLoad.scala 222:16:@3021.4]
    end
    if(tensorFile_13_0__T_6107_en & tensorFile_13_0__T_6107_mask) begin
      tensorFile_13_0[tensorFile_13_0__T_6107_addr] <= tensorFile_13_0__T_6107_data; // @[TensorLoad.scala 222:16:@3022.4]
    end
    if(tensorFile_13_1__T_6107_en & tensorFile_13_1__T_6107_mask) begin
      tensorFile_13_1[tensorFile_13_1__T_6107_addr] <= tensorFile_13_1__T_6107_data; // @[TensorLoad.scala 222:16:@3022.4]
    end
    if(tensorFile_14_0__T_6194_en & tensorFile_14_0__T_6194_mask) begin
      tensorFile_14_0[tensorFile_14_0__T_6194_addr] <= tensorFile_14_0__T_6194_data; // @[TensorLoad.scala 222:16:@3023.4]
    end
    if(tensorFile_14_1__T_6194_en & tensorFile_14_1__T_6194_mask) begin
      tensorFile_14_1[tensorFile_14_1__T_6194_addr] <= tensorFile_14_1__T_6194_data; // @[TensorLoad.scala 222:16:@3023.4]
    end
    if(tensorFile_15_0__T_6281_en & tensorFile_15_0__T_6281_mask) begin
      tensorFile_15_0[tensorFile_15_0__T_6281_addr] <= tensorFile_15_0__T_6281_data; // @[TensorLoad.scala 222:16:@3024.4]
    end
    if(tensorFile_15_1__T_6281_en & tensorFile_15_1__T_6281_mask) begin
      tensorFile_15_1[tensorFile_15_1__T_6281_addr] <= tensorFile_15_1__T_6281_data; // @[TensorLoad.scala 222:16:@3024.4]
    end
    if (reset) begin
      dataCtrlDone <= 1'h0;
    end else begin
      if (_T_4420) begin
        dataCtrlDone <= 1'h0;
      end else begin
        if (_T_4428) begin
          dataCtrlDone <= 1'h1;
        end
      end
    end
    if (_T_4492) begin
      tag <= 1'h0;
    end else begin
      if (_T_4495) begin
        tag <= _T_4498;
      end
    end
    if (_T_4506) begin
      set <= 4'h0;
    end else begin
      if (_T_4512) begin
        set <= _T_4515;
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_4394) begin
        if (io_start) begin
          if (_T_4396) begin
            state <= 3'h1;
          end else begin
            if (_T_4398) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end
      end else begin
        if (_T_4399) begin
          if (yPadCtrl0_io_done) begin
            if (_T_4398) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end else begin
          if (_T_4402) begin
            if (xPadCtrl0_io_done) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_4403) begin
              if (io_vme_rd_cmd_ready) begin
                state <= 3'h4;
              end
            end else begin
              if (_T_4404) begin
                if (io_vme_rd_data_valid) begin
                  if (dataCtrl_io_done) begin
                    if (_T_4406) begin
                      state <= 3'h5;
                    end else begin
                      if (_T_4408) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end
                  end else begin
                    if (dataCtrl_io_stride) begin
                      if (_T_4406) begin
                        state <= 3'h5;
                      end else begin
                        if (_T_4398) begin
                          state <= 3'h2;
                        end else begin
                          state <= 3'h3;
                        end
                      end
                    end else begin
                      if (dataCtrl_io_split) begin
                        state <= 3'h3;
                      end
                    end
                  end
                end
              end else begin
                if (_T_4413) begin
                  if (xPadCtrl1_io_done) begin
                    if (dataCtrlDone) begin
                      if (_T_4408) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end else begin
                      if (_T_4398) begin
                        state <= 3'h2;
                      end else begin
                        state <= 3'h3;
                      end
                    end
                  end
                end else begin
                  if (_T_4418) begin
                    if (_T_4419) begin
                      state <= 3'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    waddr_cur <= _GEN_37[9:0];
    waddr_nxt <= _GEN_38[9:0];
    rvalid <= io_tensor_rd_idx_valid;
    if (_GEN_216) begin
      tensorFile_0_0_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_0_1_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_1_0_rdata_1_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_1_1_rdata_1_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_2_0_rdata_2_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_2_1_rdata_2_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_3_0_rdata_3_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_3_1_rdata_3_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_4_0_rdata_4_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_4_1_rdata_4_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_5_0_rdata_5_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_5_1_rdata_5_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_6_0_rdata_6_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_6_1_rdata_6_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_7_0_rdata_7_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_7_1_rdata_7_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_8_0_rdata_8_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_8_1_rdata_8_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_9_0_rdata_9_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_9_1_rdata_9_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_10_0_rdata_10_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_10_1_rdata_10_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_11_0_rdata_11_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_11_1_rdata_11_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_12_0_rdata_12_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_12_1_rdata_12_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_13_0_rdata_13_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_13_1_rdata_13_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_14_0_rdata_14_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_14_1_rdata_14_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_15_0_rdata_15_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_15_1_rdata_15_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
  end
endmodule
module Load( // @[:@4857.2]
  input          clock, // @[:@4858.4]
  input          reset, // @[:@4859.4]
  input          io_i_post, // @[:@4860.4]
  output         io_o_post, // @[:@4860.4]
  output         io_inst_ready, // @[:@4860.4]
  input          io_inst_valid, // @[:@4860.4]
  input  [127:0] io_inst_bits, // @[:@4860.4]
  input  [31:0]  io_inp_baddr, // @[:@4860.4]
  input  [31:0]  io_wgt_baddr, // @[:@4860.4]
  input          io_vme_rd_0_cmd_ready, // @[:@4860.4]
  output         io_vme_rd_0_cmd_valid, // @[:@4860.4]
  output [31:0]  io_vme_rd_0_cmd_bits_addr, // @[:@4860.4]
  output [7:0]   io_vme_rd_0_cmd_bits_len, // @[:@4860.4]
  output         io_vme_rd_0_data_ready, // @[:@4860.4]
  input          io_vme_rd_0_data_valid, // @[:@4860.4]
  input  [63:0]  io_vme_rd_0_data_bits, // @[:@4860.4]
  input          io_vme_rd_1_cmd_ready, // @[:@4860.4]
  output         io_vme_rd_1_cmd_valid, // @[:@4860.4]
  output [31:0]  io_vme_rd_1_cmd_bits_addr, // @[:@4860.4]
  output [7:0]   io_vme_rd_1_cmd_bits_len, // @[:@4860.4]
  output         io_vme_rd_1_data_ready, // @[:@4860.4]
  input          io_vme_rd_1_data_valid, // @[:@4860.4]
  input  [63:0]  io_vme_rd_1_data_bits, // @[:@4860.4]
  input          io_inp_rd_idx_valid, // @[:@4860.4]
  input  [10:0]  io_inp_rd_idx_bits, // @[:@4860.4]
  output         io_inp_rd_data_valid, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_0, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_1, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_2, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_3, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_4, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_5, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_6, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_7, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_8, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_9, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_10, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_11, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_12, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_13, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_14, // @[:@4860.4]
  output [7:0]   io_inp_rd_data_bits_0_15, // @[:@4860.4]
  input          io_wgt_rd_idx_valid, // @[:@4860.4]
  input  [9:0]   io_wgt_rd_idx_bits, // @[:@4860.4]
  output         io_wgt_rd_data_valid, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_0_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_1_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_2_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_3_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_4_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_5_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_6_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_7_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_8_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_9_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_10_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_11_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_12_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_13_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_14_15, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_0, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_1, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_2, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_3, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_4, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_5, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_6, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_7, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_8, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_9, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_10, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_11, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_12, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_13, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_14, // @[:@4860.4]
  output [7:0]   io_wgt_rd_data_bits_15_15 // @[:@4860.4]
);
  wire  s_clock; // @[Load.scala 49:17:@4863.4]
  wire  s_reset; // @[Load.scala 49:17:@4863.4]
  wire  s_io_spost; // @[Load.scala 49:17:@4863.4]
  wire  s_io_swait; // @[Load.scala 49:17:@4863.4]
  wire  s_io_sready; // @[Load.scala 49:17:@4863.4]
  wire  inst_q_clock; // @[Load.scala 50:22:@4866.4]
  wire  inst_q_reset; // @[Load.scala 50:22:@4866.4]
  wire  inst_q_io_enq_ready; // @[Load.scala 50:22:@4866.4]
  wire  inst_q_io_enq_valid; // @[Load.scala 50:22:@4866.4]
  wire [127:0] inst_q_io_enq_bits; // @[Load.scala 50:22:@4866.4]
  wire  inst_q_io_deq_ready; // @[Load.scala 50:22:@4866.4]
  wire  inst_q_io_deq_valid; // @[Load.scala 50:22:@4866.4]
  wire [127:0] inst_q_io_deq_bits; // @[Load.scala 50:22:@4866.4]
  wire [127:0] dec_io_inst; // @[Load.scala 52:19:@4869.4]
  wire  dec_io_push_next; // @[Load.scala 52:19:@4869.4]
  wire  dec_io_pop_next; // @[Load.scala 52:19:@4869.4]
  wire  dec_io_isInput; // @[Load.scala 52:19:@4869.4]
  wire  dec_io_isWeight; // @[Load.scala 52:19:@4869.4]
  wire  dec_io_isSync; // @[Load.scala 52:19:@4869.4]
  wire  tensorLoad_0_clock; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_0_reset; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_0_io_start; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_0_io_done; // @[Load.scala 58:32:@4873.4]
  wire [127:0] tensorLoad_0_io_inst; // @[Load.scala 58:32:@4873.4]
  wire [31:0] tensorLoad_0_io_baddr; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_0_io_vme_rd_cmd_ready; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_0_io_vme_rd_cmd_valid; // @[Load.scala 58:32:@4873.4]
  wire [31:0] tensorLoad_0_io_vme_rd_cmd_bits_addr; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_vme_rd_cmd_bits_len; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_0_io_vme_rd_data_ready; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_0_io_vme_rd_data_valid; // @[Load.scala 58:32:@4873.4]
  wire [63:0] tensorLoad_0_io_vme_rd_data_bits; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_0_io_tensor_rd_idx_valid; // @[Load.scala 58:32:@4873.4]
  wire [10:0] tensorLoad_0_io_tensor_rd_idx_bits; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_0_io_tensor_rd_data_valid; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_0; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_1; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_2; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_3; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_4; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_5; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_6; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_7; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_8; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_9; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_10; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_11; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_12; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_13; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_14; // @[Load.scala 58:32:@4873.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_15; // @[Load.scala 58:32:@4873.4]
  wire  tensorLoad_1_clock; // @[Load.scala 58:32:@4876.4]
  wire  tensorLoad_1_reset; // @[Load.scala 58:32:@4876.4]
  wire  tensorLoad_1_io_start; // @[Load.scala 58:32:@4876.4]
  wire  tensorLoad_1_io_done; // @[Load.scala 58:32:@4876.4]
  wire [127:0] tensorLoad_1_io_inst; // @[Load.scala 58:32:@4876.4]
  wire [31:0] tensorLoad_1_io_baddr; // @[Load.scala 58:32:@4876.4]
  wire  tensorLoad_1_io_vme_rd_cmd_ready; // @[Load.scala 58:32:@4876.4]
  wire  tensorLoad_1_io_vme_rd_cmd_valid; // @[Load.scala 58:32:@4876.4]
  wire [31:0] tensorLoad_1_io_vme_rd_cmd_bits_addr; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_vme_rd_cmd_bits_len; // @[Load.scala 58:32:@4876.4]
  wire  tensorLoad_1_io_vme_rd_data_ready; // @[Load.scala 58:32:@4876.4]
  wire  tensorLoad_1_io_vme_rd_data_valid; // @[Load.scala 58:32:@4876.4]
  wire [63:0] tensorLoad_1_io_vme_rd_data_bits; // @[Load.scala 58:32:@4876.4]
  wire  tensorLoad_1_io_tensor_rd_idx_valid; // @[Load.scala 58:32:@4876.4]
  wire [9:0] tensorLoad_1_io_tensor_rd_idx_bits; // @[Load.scala 58:32:@4876.4]
  wire  tensorLoad_1_io_tensor_rd_data_valid; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_15; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_0; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_1; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_2; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_3; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_4; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_5; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_6; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_7; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_8; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_9; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_10; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_11; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_12; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_13; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_14; // @[Load.scala 58:32:@4876.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_15; // @[Load.scala 58:32:@4876.4]
  reg [1:0] state; // @[Load.scala 47:22:@4862.4]
  reg [31:0] _RAND_0;
  wire  _T_4999; // @[Load.scala 60:40:@4879.4]
  wire  start; // @[Load.scala 60:35:@4880.4]
  wire  done; // @[Load.scala 61:17:@4881.4]
  wire  _T_5000; // @[Conditional.scala 37:30:@4882.4]
  wire  _T_5001; // @[Load.scala 69:35:@4889.10]
  wire [1:0] _GEN_0; // @[Load.scala 69:55:@4890.10]
  wire [1:0] _GEN_1; // @[Load.scala 67:29:@4885.8]
  wire [1:0] _GEN_2; // @[Load.scala 66:19:@4884.6]
  wire  _T_5002; // @[Conditional.scala 37:30:@4896.6]
  wire  _T_5003; // @[Conditional.scala 37:30:@4901.8]
  wire [1:0] _GEN_3; // @[Load.scala 78:18:@4903.10]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@4902.8]
  wire [1:0] _GEN_5; // @[Conditional.scala 39:67:@4897.6]
  wire [1:0] _GEN_6; // @[Conditional.scala 40:58:@4883.4]
  wire  _T_5004; // @[Load.scala 86:33:@4910.4]
  wire  _T_5005; // @[Load.scala 86:42:@4911.4]
  wire  _T_5006; // @[Load.scala 86:59:@4912.4]
  wire  _T_5007; // @[Load.scala 86:50:@4913.4]
  wire  _T_5008; // @[Load.scala 94:37:@4915.4]
  wire  _T_5009; // @[Load.scala 94:47:@4916.4]
  Semaphore s ( // @[Load.scala 49:17:@4863.4]
    .clock(s_clock),
    .reset(s_reset),
    .io_spost(s_io_spost),
    .io_swait(s_io_swait),
    .io_sready(s_io_sready)
  );
  Queue_1 inst_q ( // @[Load.scala 50:22:@4866.4]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits)
  );
  LoadDecode dec ( // @[Load.scala 52:19:@4869.4]
    .io_inst(dec_io_inst),
    .io_push_next(dec_io_push_next),
    .io_pop_next(dec_io_pop_next),
    .io_isInput(dec_io_isInput),
    .io_isWeight(dec_io_isWeight),
    .io_isSync(dec_io_isSync)
  );
  TensorLoad tensorLoad_0 ( // @[Load.scala 58:32:@4873.4]
    .clock(tensorLoad_0_clock),
    .reset(tensorLoad_0_reset),
    .io_start(tensorLoad_0_io_start),
    .io_done(tensorLoad_0_io_done),
    .io_inst(tensorLoad_0_io_inst),
    .io_baddr(tensorLoad_0_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_0_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_0_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_0_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_0_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(tensorLoad_0_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorLoad_0_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(tensorLoad_0_io_vme_rd_data_bits),
    .io_tensor_rd_idx_valid(tensorLoad_0_io_tensor_rd_idx_valid),
    .io_tensor_rd_idx_bits(tensorLoad_0_io_tensor_rd_idx_bits),
    .io_tensor_rd_data_valid(tensorLoad_0_io_tensor_rd_data_valid),
    .io_tensor_rd_data_bits_0_0(tensorLoad_0_io_tensor_rd_data_bits_0_0),
    .io_tensor_rd_data_bits_0_1(tensorLoad_0_io_tensor_rd_data_bits_0_1),
    .io_tensor_rd_data_bits_0_2(tensorLoad_0_io_tensor_rd_data_bits_0_2),
    .io_tensor_rd_data_bits_0_3(tensorLoad_0_io_tensor_rd_data_bits_0_3),
    .io_tensor_rd_data_bits_0_4(tensorLoad_0_io_tensor_rd_data_bits_0_4),
    .io_tensor_rd_data_bits_0_5(tensorLoad_0_io_tensor_rd_data_bits_0_5),
    .io_tensor_rd_data_bits_0_6(tensorLoad_0_io_tensor_rd_data_bits_0_6),
    .io_tensor_rd_data_bits_0_7(tensorLoad_0_io_tensor_rd_data_bits_0_7),
    .io_tensor_rd_data_bits_0_8(tensorLoad_0_io_tensor_rd_data_bits_0_8),
    .io_tensor_rd_data_bits_0_9(tensorLoad_0_io_tensor_rd_data_bits_0_9),
    .io_tensor_rd_data_bits_0_10(tensorLoad_0_io_tensor_rd_data_bits_0_10),
    .io_tensor_rd_data_bits_0_11(tensorLoad_0_io_tensor_rd_data_bits_0_11),
    .io_tensor_rd_data_bits_0_12(tensorLoad_0_io_tensor_rd_data_bits_0_12),
    .io_tensor_rd_data_bits_0_13(tensorLoad_0_io_tensor_rd_data_bits_0_13),
    .io_tensor_rd_data_bits_0_14(tensorLoad_0_io_tensor_rd_data_bits_0_14),
    .io_tensor_rd_data_bits_0_15(tensorLoad_0_io_tensor_rd_data_bits_0_15)
  );
  TensorLoad_1 tensorLoad_1 ( // @[Load.scala 58:32:@4876.4]
    .clock(tensorLoad_1_clock),
    .reset(tensorLoad_1_reset),
    .io_start(tensorLoad_1_io_start),
    .io_done(tensorLoad_1_io_done),
    .io_inst(tensorLoad_1_io_inst),
    .io_baddr(tensorLoad_1_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_1_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_1_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_1_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_1_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(tensorLoad_1_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorLoad_1_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(tensorLoad_1_io_vme_rd_data_bits),
    .io_tensor_rd_idx_valid(tensorLoad_1_io_tensor_rd_idx_valid),
    .io_tensor_rd_idx_bits(tensorLoad_1_io_tensor_rd_idx_bits),
    .io_tensor_rd_data_valid(tensorLoad_1_io_tensor_rd_data_valid),
    .io_tensor_rd_data_bits_0_0(tensorLoad_1_io_tensor_rd_data_bits_0_0),
    .io_tensor_rd_data_bits_0_1(tensorLoad_1_io_tensor_rd_data_bits_0_1),
    .io_tensor_rd_data_bits_0_2(tensorLoad_1_io_tensor_rd_data_bits_0_2),
    .io_tensor_rd_data_bits_0_3(tensorLoad_1_io_tensor_rd_data_bits_0_3),
    .io_tensor_rd_data_bits_0_4(tensorLoad_1_io_tensor_rd_data_bits_0_4),
    .io_tensor_rd_data_bits_0_5(tensorLoad_1_io_tensor_rd_data_bits_0_5),
    .io_tensor_rd_data_bits_0_6(tensorLoad_1_io_tensor_rd_data_bits_0_6),
    .io_tensor_rd_data_bits_0_7(tensorLoad_1_io_tensor_rd_data_bits_0_7),
    .io_tensor_rd_data_bits_0_8(tensorLoad_1_io_tensor_rd_data_bits_0_8),
    .io_tensor_rd_data_bits_0_9(tensorLoad_1_io_tensor_rd_data_bits_0_9),
    .io_tensor_rd_data_bits_0_10(tensorLoad_1_io_tensor_rd_data_bits_0_10),
    .io_tensor_rd_data_bits_0_11(tensorLoad_1_io_tensor_rd_data_bits_0_11),
    .io_tensor_rd_data_bits_0_12(tensorLoad_1_io_tensor_rd_data_bits_0_12),
    .io_tensor_rd_data_bits_0_13(tensorLoad_1_io_tensor_rd_data_bits_0_13),
    .io_tensor_rd_data_bits_0_14(tensorLoad_1_io_tensor_rd_data_bits_0_14),
    .io_tensor_rd_data_bits_0_15(tensorLoad_1_io_tensor_rd_data_bits_0_15),
    .io_tensor_rd_data_bits_1_0(tensorLoad_1_io_tensor_rd_data_bits_1_0),
    .io_tensor_rd_data_bits_1_1(tensorLoad_1_io_tensor_rd_data_bits_1_1),
    .io_tensor_rd_data_bits_1_2(tensorLoad_1_io_tensor_rd_data_bits_1_2),
    .io_tensor_rd_data_bits_1_3(tensorLoad_1_io_tensor_rd_data_bits_1_3),
    .io_tensor_rd_data_bits_1_4(tensorLoad_1_io_tensor_rd_data_bits_1_4),
    .io_tensor_rd_data_bits_1_5(tensorLoad_1_io_tensor_rd_data_bits_1_5),
    .io_tensor_rd_data_bits_1_6(tensorLoad_1_io_tensor_rd_data_bits_1_6),
    .io_tensor_rd_data_bits_1_7(tensorLoad_1_io_tensor_rd_data_bits_1_7),
    .io_tensor_rd_data_bits_1_8(tensorLoad_1_io_tensor_rd_data_bits_1_8),
    .io_tensor_rd_data_bits_1_9(tensorLoad_1_io_tensor_rd_data_bits_1_9),
    .io_tensor_rd_data_bits_1_10(tensorLoad_1_io_tensor_rd_data_bits_1_10),
    .io_tensor_rd_data_bits_1_11(tensorLoad_1_io_tensor_rd_data_bits_1_11),
    .io_tensor_rd_data_bits_1_12(tensorLoad_1_io_tensor_rd_data_bits_1_12),
    .io_tensor_rd_data_bits_1_13(tensorLoad_1_io_tensor_rd_data_bits_1_13),
    .io_tensor_rd_data_bits_1_14(tensorLoad_1_io_tensor_rd_data_bits_1_14),
    .io_tensor_rd_data_bits_1_15(tensorLoad_1_io_tensor_rd_data_bits_1_15),
    .io_tensor_rd_data_bits_2_0(tensorLoad_1_io_tensor_rd_data_bits_2_0),
    .io_tensor_rd_data_bits_2_1(tensorLoad_1_io_tensor_rd_data_bits_2_1),
    .io_tensor_rd_data_bits_2_2(tensorLoad_1_io_tensor_rd_data_bits_2_2),
    .io_tensor_rd_data_bits_2_3(tensorLoad_1_io_tensor_rd_data_bits_2_3),
    .io_tensor_rd_data_bits_2_4(tensorLoad_1_io_tensor_rd_data_bits_2_4),
    .io_tensor_rd_data_bits_2_5(tensorLoad_1_io_tensor_rd_data_bits_2_5),
    .io_tensor_rd_data_bits_2_6(tensorLoad_1_io_tensor_rd_data_bits_2_6),
    .io_tensor_rd_data_bits_2_7(tensorLoad_1_io_tensor_rd_data_bits_2_7),
    .io_tensor_rd_data_bits_2_8(tensorLoad_1_io_tensor_rd_data_bits_2_8),
    .io_tensor_rd_data_bits_2_9(tensorLoad_1_io_tensor_rd_data_bits_2_9),
    .io_tensor_rd_data_bits_2_10(tensorLoad_1_io_tensor_rd_data_bits_2_10),
    .io_tensor_rd_data_bits_2_11(tensorLoad_1_io_tensor_rd_data_bits_2_11),
    .io_tensor_rd_data_bits_2_12(tensorLoad_1_io_tensor_rd_data_bits_2_12),
    .io_tensor_rd_data_bits_2_13(tensorLoad_1_io_tensor_rd_data_bits_2_13),
    .io_tensor_rd_data_bits_2_14(tensorLoad_1_io_tensor_rd_data_bits_2_14),
    .io_tensor_rd_data_bits_2_15(tensorLoad_1_io_tensor_rd_data_bits_2_15),
    .io_tensor_rd_data_bits_3_0(tensorLoad_1_io_tensor_rd_data_bits_3_0),
    .io_tensor_rd_data_bits_3_1(tensorLoad_1_io_tensor_rd_data_bits_3_1),
    .io_tensor_rd_data_bits_3_2(tensorLoad_1_io_tensor_rd_data_bits_3_2),
    .io_tensor_rd_data_bits_3_3(tensorLoad_1_io_tensor_rd_data_bits_3_3),
    .io_tensor_rd_data_bits_3_4(tensorLoad_1_io_tensor_rd_data_bits_3_4),
    .io_tensor_rd_data_bits_3_5(tensorLoad_1_io_tensor_rd_data_bits_3_5),
    .io_tensor_rd_data_bits_3_6(tensorLoad_1_io_tensor_rd_data_bits_3_6),
    .io_tensor_rd_data_bits_3_7(tensorLoad_1_io_tensor_rd_data_bits_3_7),
    .io_tensor_rd_data_bits_3_8(tensorLoad_1_io_tensor_rd_data_bits_3_8),
    .io_tensor_rd_data_bits_3_9(tensorLoad_1_io_tensor_rd_data_bits_3_9),
    .io_tensor_rd_data_bits_3_10(tensorLoad_1_io_tensor_rd_data_bits_3_10),
    .io_tensor_rd_data_bits_3_11(tensorLoad_1_io_tensor_rd_data_bits_3_11),
    .io_tensor_rd_data_bits_3_12(tensorLoad_1_io_tensor_rd_data_bits_3_12),
    .io_tensor_rd_data_bits_3_13(tensorLoad_1_io_tensor_rd_data_bits_3_13),
    .io_tensor_rd_data_bits_3_14(tensorLoad_1_io_tensor_rd_data_bits_3_14),
    .io_tensor_rd_data_bits_3_15(tensorLoad_1_io_tensor_rd_data_bits_3_15),
    .io_tensor_rd_data_bits_4_0(tensorLoad_1_io_tensor_rd_data_bits_4_0),
    .io_tensor_rd_data_bits_4_1(tensorLoad_1_io_tensor_rd_data_bits_4_1),
    .io_tensor_rd_data_bits_4_2(tensorLoad_1_io_tensor_rd_data_bits_4_2),
    .io_tensor_rd_data_bits_4_3(tensorLoad_1_io_tensor_rd_data_bits_4_3),
    .io_tensor_rd_data_bits_4_4(tensorLoad_1_io_tensor_rd_data_bits_4_4),
    .io_tensor_rd_data_bits_4_5(tensorLoad_1_io_tensor_rd_data_bits_4_5),
    .io_tensor_rd_data_bits_4_6(tensorLoad_1_io_tensor_rd_data_bits_4_6),
    .io_tensor_rd_data_bits_4_7(tensorLoad_1_io_tensor_rd_data_bits_4_7),
    .io_tensor_rd_data_bits_4_8(tensorLoad_1_io_tensor_rd_data_bits_4_8),
    .io_tensor_rd_data_bits_4_9(tensorLoad_1_io_tensor_rd_data_bits_4_9),
    .io_tensor_rd_data_bits_4_10(tensorLoad_1_io_tensor_rd_data_bits_4_10),
    .io_tensor_rd_data_bits_4_11(tensorLoad_1_io_tensor_rd_data_bits_4_11),
    .io_tensor_rd_data_bits_4_12(tensorLoad_1_io_tensor_rd_data_bits_4_12),
    .io_tensor_rd_data_bits_4_13(tensorLoad_1_io_tensor_rd_data_bits_4_13),
    .io_tensor_rd_data_bits_4_14(tensorLoad_1_io_tensor_rd_data_bits_4_14),
    .io_tensor_rd_data_bits_4_15(tensorLoad_1_io_tensor_rd_data_bits_4_15),
    .io_tensor_rd_data_bits_5_0(tensorLoad_1_io_tensor_rd_data_bits_5_0),
    .io_tensor_rd_data_bits_5_1(tensorLoad_1_io_tensor_rd_data_bits_5_1),
    .io_tensor_rd_data_bits_5_2(tensorLoad_1_io_tensor_rd_data_bits_5_2),
    .io_tensor_rd_data_bits_5_3(tensorLoad_1_io_tensor_rd_data_bits_5_3),
    .io_tensor_rd_data_bits_5_4(tensorLoad_1_io_tensor_rd_data_bits_5_4),
    .io_tensor_rd_data_bits_5_5(tensorLoad_1_io_tensor_rd_data_bits_5_5),
    .io_tensor_rd_data_bits_5_6(tensorLoad_1_io_tensor_rd_data_bits_5_6),
    .io_tensor_rd_data_bits_5_7(tensorLoad_1_io_tensor_rd_data_bits_5_7),
    .io_tensor_rd_data_bits_5_8(tensorLoad_1_io_tensor_rd_data_bits_5_8),
    .io_tensor_rd_data_bits_5_9(tensorLoad_1_io_tensor_rd_data_bits_5_9),
    .io_tensor_rd_data_bits_5_10(tensorLoad_1_io_tensor_rd_data_bits_5_10),
    .io_tensor_rd_data_bits_5_11(tensorLoad_1_io_tensor_rd_data_bits_5_11),
    .io_tensor_rd_data_bits_5_12(tensorLoad_1_io_tensor_rd_data_bits_5_12),
    .io_tensor_rd_data_bits_5_13(tensorLoad_1_io_tensor_rd_data_bits_5_13),
    .io_tensor_rd_data_bits_5_14(tensorLoad_1_io_tensor_rd_data_bits_5_14),
    .io_tensor_rd_data_bits_5_15(tensorLoad_1_io_tensor_rd_data_bits_5_15),
    .io_tensor_rd_data_bits_6_0(tensorLoad_1_io_tensor_rd_data_bits_6_0),
    .io_tensor_rd_data_bits_6_1(tensorLoad_1_io_tensor_rd_data_bits_6_1),
    .io_tensor_rd_data_bits_6_2(tensorLoad_1_io_tensor_rd_data_bits_6_2),
    .io_tensor_rd_data_bits_6_3(tensorLoad_1_io_tensor_rd_data_bits_6_3),
    .io_tensor_rd_data_bits_6_4(tensorLoad_1_io_tensor_rd_data_bits_6_4),
    .io_tensor_rd_data_bits_6_5(tensorLoad_1_io_tensor_rd_data_bits_6_5),
    .io_tensor_rd_data_bits_6_6(tensorLoad_1_io_tensor_rd_data_bits_6_6),
    .io_tensor_rd_data_bits_6_7(tensorLoad_1_io_tensor_rd_data_bits_6_7),
    .io_tensor_rd_data_bits_6_8(tensorLoad_1_io_tensor_rd_data_bits_6_8),
    .io_tensor_rd_data_bits_6_9(tensorLoad_1_io_tensor_rd_data_bits_6_9),
    .io_tensor_rd_data_bits_6_10(tensorLoad_1_io_tensor_rd_data_bits_6_10),
    .io_tensor_rd_data_bits_6_11(tensorLoad_1_io_tensor_rd_data_bits_6_11),
    .io_tensor_rd_data_bits_6_12(tensorLoad_1_io_tensor_rd_data_bits_6_12),
    .io_tensor_rd_data_bits_6_13(tensorLoad_1_io_tensor_rd_data_bits_6_13),
    .io_tensor_rd_data_bits_6_14(tensorLoad_1_io_tensor_rd_data_bits_6_14),
    .io_tensor_rd_data_bits_6_15(tensorLoad_1_io_tensor_rd_data_bits_6_15),
    .io_tensor_rd_data_bits_7_0(tensorLoad_1_io_tensor_rd_data_bits_7_0),
    .io_tensor_rd_data_bits_7_1(tensorLoad_1_io_tensor_rd_data_bits_7_1),
    .io_tensor_rd_data_bits_7_2(tensorLoad_1_io_tensor_rd_data_bits_7_2),
    .io_tensor_rd_data_bits_7_3(tensorLoad_1_io_tensor_rd_data_bits_7_3),
    .io_tensor_rd_data_bits_7_4(tensorLoad_1_io_tensor_rd_data_bits_7_4),
    .io_tensor_rd_data_bits_7_5(tensorLoad_1_io_tensor_rd_data_bits_7_5),
    .io_tensor_rd_data_bits_7_6(tensorLoad_1_io_tensor_rd_data_bits_7_6),
    .io_tensor_rd_data_bits_7_7(tensorLoad_1_io_tensor_rd_data_bits_7_7),
    .io_tensor_rd_data_bits_7_8(tensorLoad_1_io_tensor_rd_data_bits_7_8),
    .io_tensor_rd_data_bits_7_9(tensorLoad_1_io_tensor_rd_data_bits_7_9),
    .io_tensor_rd_data_bits_7_10(tensorLoad_1_io_tensor_rd_data_bits_7_10),
    .io_tensor_rd_data_bits_7_11(tensorLoad_1_io_tensor_rd_data_bits_7_11),
    .io_tensor_rd_data_bits_7_12(tensorLoad_1_io_tensor_rd_data_bits_7_12),
    .io_tensor_rd_data_bits_7_13(tensorLoad_1_io_tensor_rd_data_bits_7_13),
    .io_tensor_rd_data_bits_7_14(tensorLoad_1_io_tensor_rd_data_bits_7_14),
    .io_tensor_rd_data_bits_7_15(tensorLoad_1_io_tensor_rd_data_bits_7_15),
    .io_tensor_rd_data_bits_8_0(tensorLoad_1_io_tensor_rd_data_bits_8_0),
    .io_tensor_rd_data_bits_8_1(tensorLoad_1_io_tensor_rd_data_bits_8_1),
    .io_tensor_rd_data_bits_8_2(tensorLoad_1_io_tensor_rd_data_bits_8_2),
    .io_tensor_rd_data_bits_8_3(tensorLoad_1_io_tensor_rd_data_bits_8_3),
    .io_tensor_rd_data_bits_8_4(tensorLoad_1_io_tensor_rd_data_bits_8_4),
    .io_tensor_rd_data_bits_8_5(tensorLoad_1_io_tensor_rd_data_bits_8_5),
    .io_tensor_rd_data_bits_8_6(tensorLoad_1_io_tensor_rd_data_bits_8_6),
    .io_tensor_rd_data_bits_8_7(tensorLoad_1_io_tensor_rd_data_bits_8_7),
    .io_tensor_rd_data_bits_8_8(tensorLoad_1_io_tensor_rd_data_bits_8_8),
    .io_tensor_rd_data_bits_8_9(tensorLoad_1_io_tensor_rd_data_bits_8_9),
    .io_tensor_rd_data_bits_8_10(tensorLoad_1_io_tensor_rd_data_bits_8_10),
    .io_tensor_rd_data_bits_8_11(tensorLoad_1_io_tensor_rd_data_bits_8_11),
    .io_tensor_rd_data_bits_8_12(tensorLoad_1_io_tensor_rd_data_bits_8_12),
    .io_tensor_rd_data_bits_8_13(tensorLoad_1_io_tensor_rd_data_bits_8_13),
    .io_tensor_rd_data_bits_8_14(tensorLoad_1_io_tensor_rd_data_bits_8_14),
    .io_tensor_rd_data_bits_8_15(tensorLoad_1_io_tensor_rd_data_bits_8_15),
    .io_tensor_rd_data_bits_9_0(tensorLoad_1_io_tensor_rd_data_bits_9_0),
    .io_tensor_rd_data_bits_9_1(tensorLoad_1_io_tensor_rd_data_bits_9_1),
    .io_tensor_rd_data_bits_9_2(tensorLoad_1_io_tensor_rd_data_bits_9_2),
    .io_tensor_rd_data_bits_9_3(tensorLoad_1_io_tensor_rd_data_bits_9_3),
    .io_tensor_rd_data_bits_9_4(tensorLoad_1_io_tensor_rd_data_bits_9_4),
    .io_tensor_rd_data_bits_9_5(tensorLoad_1_io_tensor_rd_data_bits_9_5),
    .io_tensor_rd_data_bits_9_6(tensorLoad_1_io_tensor_rd_data_bits_9_6),
    .io_tensor_rd_data_bits_9_7(tensorLoad_1_io_tensor_rd_data_bits_9_7),
    .io_tensor_rd_data_bits_9_8(tensorLoad_1_io_tensor_rd_data_bits_9_8),
    .io_tensor_rd_data_bits_9_9(tensorLoad_1_io_tensor_rd_data_bits_9_9),
    .io_tensor_rd_data_bits_9_10(tensorLoad_1_io_tensor_rd_data_bits_9_10),
    .io_tensor_rd_data_bits_9_11(tensorLoad_1_io_tensor_rd_data_bits_9_11),
    .io_tensor_rd_data_bits_9_12(tensorLoad_1_io_tensor_rd_data_bits_9_12),
    .io_tensor_rd_data_bits_9_13(tensorLoad_1_io_tensor_rd_data_bits_9_13),
    .io_tensor_rd_data_bits_9_14(tensorLoad_1_io_tensor_rd_data_bits_9_14),
    .io_tensor_rd_data_bits_9_15(tensorLoad_1_io_tensor_rd_data_bits_9_15),
    .io_tensor_rd_data_bits_10_0(tensorLoad_1_io_tensor_rd_data_bits_10_0),
    .io_tensor_rd_data_bits_10_1(tensorLoad_1_io_tensor_rd_data_bits_10_1),
    .io_tensor_rd_data_bits_10_2(tensorLoad_1_io_tensor_rd_data_bits_10_2),
    .io_tensor_rd_data_bits_10_3(tensorLoad_1_io_tensor_rd_data_bits_10_3),
    .io_tensor_rd_data_bits_10_4(tensorLoad_1_io_tensor_rd_data_bits_10_4),
    .io_tensor_rd_data_bits_10_5(tensorLoad_1_io_tensor_rd_data_bits_10_5),
    .io_tensor_rd_data_bits_10_6(tensorLoad_1_io_tensor_rd_data_bits_10_6),
    .io_tensor_rd_data_bits_10_7(tensorLoad_1_io_tensor_rd_data_bits_10_7),
    .io_tensor_rd_data_bits_10_8(tensorLoad_1_io_tensor_rd_data_bits_10_8),
    .io_tensor_rd_data_bits_10_9(tensorLoad_1_io_tensor_rd_data_bits_10_9),
    .io_tensor_rd_data_bits_10_10(tensorLoad_1_io_tensor_rd_data_bits_10_10),
    .io_tensor_rd_data_bits_10_11(tensorLoad_1_io_tensor_rd_data_bits_10_11),
    .io_tensor_rd_data_bits_10_12(tensorLoad_1_io_tensor_rd_data_bits_10_12),
    .io_tensor_rd_data_bits_10_13(tensorLoad_1_io_tensor_rd_data_bits_10_13),
    .io_tensor_rd_data_bits_10_14(tensorLoad_1_io_tensor_rd_data_bits_10_14),
    .io_tensor_rd_data_bits_10_15(tensorLoad_1_io_tensor_rd_data_bits_10_15),
    .io_tensor_rd_data_bits_11_0(tensorLoad_1_io_tensor_rd_data_bits_11_0),
    .io_tensor_rd_data_bits_11_1(tensorLoad_1_io_tensor_rd_data_bits_11_1),
    .io_tensor_rd_data_bits_11_2(tensorLoad_1_io_tensor_rd_data_bits_11_2),
    .io_tensor_rd_data_bits_11_3(tensorLoad_1_io_tensor_rd_data_bits_11_3),
    .io_tensor_rd_data_bits_11_4(tensorLoad_1_io_tensor_rd_data_bits_11_4),
    .io_tensor_rd_data_bits_11_5(tensorLoad_1_io_tensor_rd_data_bits_11_5),
    .io_tensor_rd_data_bits_11_6(tensorLoad_1_io_tensor_rd_data_bits_11_6),
    .io_tensor_rd_data_bits_11_7(tensorLoad_1_io_tensor_rd_data_bits_11_7),
    .io_tensor_rd_data_bits_11_8(tensorLoad_1_io_tensor_rd_data_bits_11_8),
    .io_tensor_rd_data_bits_11_9(tensorLoad_1_io_tensor_rd_data_bits_11_9),
    .io_tensor_rd_data_bits_11_10(tensorLoad_1_io_tensor_rd_data_bits_11_10),
    .io_tensor_rd_data_bits_11_11(tensorLoad_1_io_tensor_rd_data_bits_11_11),
    .io_tensor_rd_data_bits_11_12(tensorLoad_1_io_tensor_rd_data_bits_11_12),
    .io_tensor_rd_data_bits_11_13(tensorLoad_1_io_tensor_rd_data_bits_11_13),
    .io_tensor_rd_data_bits_11_14(tensorLoad_1_io_tensor_rd_data_bits_11_14),
    .io_tensor_rd_data_bits_11_15(tensorLoad_1_io_tensor_rd_data_bits_11_15),
    .io_tensor_rd_data_bits_12_0(tensorLoad_1_io_tensor_rd_data_bits_12_0),
    .io_tensor_rd_data_bits_12_1(tensorLoad_1_io_tensor_rd_data_bits_12_1),
    .io_tensor_rd_data_bits_12_2(tensorLoad_1_io_tensor_rd_data_bits_12_2),
    .io_tensor_rd_data_bits_12_3(tensorLoad_1_io_tensor_rd_data_bits_12_3),
    .io_tensor_rd_data_bits_12_4(tensorLoad_1_io_tensor_rd_data_bits_12_4),
    .io_tensor_rd_data_bits_12_5(tensorLoad_1_io_tensor_rd_data_bits_12_5),
    .io_tensor_rd_data_bits_12_6(tensorLoad_1_io_tensor_rd_data_bits_12_6),
    .io_tensor_rd_data_bits_12_7(tensorLoad_1_io_tensor_rd_data_bits_12_7),
    .io_tensor_rd_data_bits_12_8(tensorLoad_1_io_tensor_rd_data_bits_12_8),
    .io_tensor_rd_data_bits_12_9(tensorLoad_1_io_tensor_rd_data_bits_12_9),
    .io_tensor_rd_data_bits_12_10(tensorLoad_1_io_tensor_rd_data_bits_12_10),
    .io_tensor_rd_data_bits_12_11(tensorLoad_1_io_tensor_rd_data_bits_12_11),
    .io_tensor_rd_data_bits_12_12(tensorLoad_1_io_tensor_rd_data_bits_12_12),
    .io_tensor_rd_data_bits_12_13(tensorLoad_1_io_tensor_rd_data_bits_12_13),
    .io_tensor_rd_data_bits_12_14(tensorLoad_1_io_tensor_rd_data_bits_12_14),
    .io_tensor_rd_data_bits_12_15(tensorLoad_1_io_tensor_rd_data_bits_12_15),
    .io_tensor_rd_data_bits_13_0(tensorLoad_1_io_tensor_rd_data_bits_13_0),
    .io_tensor_rd_data_bits_13_1(tensorLoad_1_io_tensor_rd_data_bits_13_1),
    .io_tensor_rd_data_bits_13_2(tensorLoad_1_io_tensor_rd_data_bits_13_2),
    .io_tensor_rd_data_bits_13_3(tensorLoad_1_io_tensor_rd_data_bits_13_3),
    .io_tensor_rd_data_bits_13_4(tensorLoad_1_io_tensor_rd_data_bits_13_4),
    .io_tensor_rd_data_bits_13_5(tensorLoad_1_io_tensor_rd_data_bits_13_5),
    .io_tensor_rd_data_bits_13_6(tensorLoad_1_io_tensor_rd_data_bits_13_6),
    .io_tensor_rd_data_bits_13_7(tensorLoad_1_io_tensor_rd_data_bits_13_7),
    .io_tensor_rd_data_bits_13_8(tensorLoad_1_io_tensor_rd_data_bits_13_8),
    .io_tensor_rd_data_bits_13_9(tensorLoad_1_io_tensor_rd_data_bits_13_9),
    .io_tensor_rd_data_bits_13_10(tensorLoad_1_io_tensor_rd_data_bits_13_10),
    .io_tensor_rd_data_bits_13_11(tensorLoad_1_io_tensor_rd_data_bits_13_11),
    .io_tensor_rd_data_bits_13_12(tensorLoad_1_io_tensor_rd_data_bits_13_12),
    .io_tensor_rd_data_bits_13_13(tensorLoad_1_io_tensor_rd_data_bits_13_13),
    .io_tensor_rd_data_bits_13_14(tensorLoad_1_io_tensor_rd_data_bits_13_14),
    .io_tensor_rd_data_bits_13_15(tensorLoad_1_io_tensor_rd_data_bits_13_15),
    .io_tensor_rd_data_bits_14_0(tensorLoad_1_io_tensor_rd_data_bits_14_0),
    .io_tensor_rd_data_bits_14_1(tensorLoad_1_io_tensor_rd_data_bits_14_1),
    .io_tensor_rd_data_bits_14_2(tensorLoad_1_io_tensor_rd_data_bits_14_2),
    .io_tensor_rd_data_bits_14_3(tensorLoad_1_io_tensor_rd_data_bits_14_3),
    .io_tensor_rd_data_bits_14_4(tensorLoad_1_io_tensor_rd_data_bits_14_4),
    .io_tensor_rd_data_bits_14_5(tensorLoad_1_io_tensor_rd_data_bits_14_5),
    .io_tensor_rd_data_bits_14_6(tensorLoad_1_io_tensor_rd_data_bits_14_6),
    .io_tensor_rd_data_bits_14_7(tensorLoad_1_io_tensor_rd_data_bits_14_7),
    .io_tensor_rd_data_bits_14_8(tensorLoad_1_io_tensor_rd_data_bits_14_8),
    .io_tensor_rd_data_bits_14_9(tensorLoad_1_io_tensor_rd_data_bits_14_9),
    .io_tensor_rd_data_bits_14_10(tensorLoad_1_io_tensor_rd_data_bits_14_10),
    .io_tensor_rd_data_bits_14_11(tensorLoad_1_io_tensor_rd_data_bits_14_11),
    .io_tensor_rd_data_bits_14_12(tensorLoad_1_io_tensor_rd_data_bits_14_12),
    .io_tensor_rd_data_bits_14_13(tensorLoad_1_io_tensor_rd_data_bits_14_13),
    .io_tensor_rd_data_bits_14_14(tensorLoad_1_io_tensor_rd_data_bits_14_14),
    .io_tensor_rd_data_bits_14_15(tensorLoad_1_io_tensor_rd_data_bits_14_15),
    .io_tensor_rd_data_bits_15_0(tensorLoad_1_io_tensor_rd_data_bits_15_0),
    .io_tensor_rd_data_bits_15_1(tensorLoad_1_io_tensor_rd_data_bits_15_1),
    .io_tensor_rd_data_bits_15_2(tensorLoad_1_io_tensor_rd_data_bits_15_2),
    .io_tensor_rd_data_bits_15_3(tensorLoad_1_io_tensor_rd_data_bits_15_3),
    .io_tensor_rd_data_bits_15_4(tensorLoad_1_io_tensor_rd_data_bits_15_4),
    .io_tensor_rd_data_bits_15_5(tensorLoad_1_io_tensor_rd_data_bits_15_5),
    .io_tensor_rd_data_bits_15_6(tensorLoad_1_io_tensor_rd_data_bits_15_6),
    .io_tensor_rd_data_bits_15_7(tensorLoad_1_io_tensor_rd_data_bits_15_7),
    .io_tensor_rd_data_bits_15_8(tensorLoad_1_io_tensor_rd_data_bits_15_8),
    .io_tensor_rd_data_bits_15_9(tensorLoad_1_io_tensor_rd_data_bits_15_9),
    .io_tensor_rd_data_bits_15_10(tensorLoad_1_io_tensor_rd_data_bits_15_10),
    .io_tensor_rd_data_bits_15_11(tensorLoad_1_io_tensor_rd_data_bits_15_11),
    .io_tensor_rd_data_bits_15_12(tensorLoad_1_io_tensor_rd_data_bits_15_12),
    .io_tensor_rd_data_bits_15_13(tensorLoad_1_io_tensor_rd_data_bits_15_13),
    .io_tensor_rd_data_bits_15_14(tensorLoad_1_io_tensor_rd_data_bits_15_14),
    .io_tensor_rd_data_bits_15_15(tensorLoad_1_io_tensor_rd_data_bits_15_15)
  );
  assign _T_4999 = dec_io_pop_next ? s_io_sready : 1'h1; // @[Load.scala 60:40:@4879.4]
  assign start = inst_q_io_deq_valid & _T_4999; // @[Load.scala 60:35:@4880.4]
  assign done = dec_io_isInput ? tensorLoad_0_io_done : tensorLoad_1_io_done; // @[Load.scala 61:17:@4881.4]
  assign _T_5000 = 2'h0 == state; // @[Conditional.scala 37:30:@4882.4]
  assign _T_5001 = dec_io_isInput | dec_io_isWeight; // @[Load.scala 69:35:@4889.10]
  assign _GEN_0 = _T_5001 ? 2'h2 : state; // @[Load.scala 69:55:@4890.10]
  assign _GEN_1 = dec_io_isSync ? 2'h1 : _GEN_0; // @[Load.scala 67:29:@4885.8]
  assign _GEN_2 = start ? _GEN_1 : state; // @[Load.scala 66:19:@4884.6]
  assign _T_5002 = 2'h1 == state; // @[Conditional.scala 37:30:@4896.6]
  assign _T_5003 = 2'h2 == state; // @[Conditional.scala 37:30:@4901.8]
  assign _GEN_3 = done ? 2'h0 : state; // @[Load.scala 78:18:@4903.10]
  assign _GEN_4 = _T_5003 ? _GEN_3 : state; // @[Conditional.scala 39:67:@4902.8]
  assign _GEN_5 = _T_5002 ? 2'h0 : _GEN_4; // @[Conditional.scala 39:67:@4897.6]
  assign _GEN_6 = _T_5000 ? _GEN_2 : _GEN_5; // @[Conditional.scala 40:58:@4883.4]
  assign _T_5004 = state == 2'h2; // @[Load.scala 86:33:@4910.4]
  assign _T_5005 = _T_5004 & done; // @[Load.scala 86:42:@4911.4]
  assign _T_5006 = state == 2'h1; // @[Load.scala 86:59:@4912.4]
  assign _T_5007 = _T_5005 | _T_5006; // @[Load.scala 86:50:@4913.4]
  assign _T_5008 = state == 2'h0; // @[Load.scala 94:37:@4915.4]
  assign _T_5009 = _T_5008 & start; // @[Load.scala 94:47:@4916.4]
  assign io_o_post = dec_io_push_next & _T_5007; // @[Load.scala 104:13:@5505.4]
  assign io_inst_ready = inst_q_io_enq_ready; // @[Load.scala 85:17:@4909.4]
  assign io_vme_rd_0_cmd_valid = tensorLoad_0_io_vme_rd_cmd_valid; // @[Load.scala 98:18:@4963.4]
  assign io_vme_rd_0_cmd_bits_addr = tensorLoad_0_io_vme_rd_cmd_bits_addr; // @[Load.scala 98:18:@4962.4]
  assign io_vme_rd_0_cmd_bits_len = tensorLoad_0_io_vme_rd_cmd_bits_len; // @[Load.scala 98:18:@4961.4]
  assign io_vme_rd_0_data_ready = tensorLoad_0_io_vme_rd_data_ready; // @[Load.scala 98:18:@4960.4]
  assign io_vme_rd_1_cmd_valid = tensorLoad_1_io_vme_rd_cmd_valid; // @[Load.scala 98:18:@5493.4]
  assign io_vme_rd_1_cmd_bits_addr = tensorLoad_1_io_vme_rd_cmd_bits_addr; // @[Load.scala 98:18:@5492.4]
  assign io_vme_rd_1_cmd_bits_len = tensorLoad_1_io_vme_rd_cmd_bits_len; // @[Load.scala 98:18:@5491.4]
  assign io_vme_rd_1_data_ready = tensorLoad_1_io_vme_rd_data_ready; // @[Load.scala 98:18:@5490.4]
  assign io_inp_rd_data_valid = tensorLoad_0_io_tensor_rd_data_valid; // @[Load.scala 97:29:@4955.4]
  assign io_inp_rd_data_bits_0_0 = tensorLoad_0_io_tensor_rd_data_bits_0_0; // @[Load.scala 97:29:@4939.4]
  assign io_inp_rd_data_bits_0_1 = tensorLoad_0_io_tensor_rd_data_bits_0_1; // @[Load.scala 97:29:@4940.4]
  assign io_inp_rd_data_bits_0_2 = tensorLoad_0_io_tensor_rd_data_bits_0_2; // @[Load.scala 97:29:@4941.4]
  assign io_inp_rd_data_bits_0_3 = tensorLoad_0_io_tensor_rd_data_bits_0_3; // @[Load.scala 97:29:@4942.4]
  assign io_inp_rd_data_bits_0_4 = tensorLoad_0_io_tensor_rd_data_bits_0_4; // @[Load.scala 97:29:@4943.4]
  assign io_inp_rd_data_bits_0_5 = tensorLoad_0_io_tensor_rd_data_bits_0_5; // @[Load.scala 97:29:@4944.4]
  assign io_inp_rd_data_bits_0_6 = tensorLoad_0_io_tensor_rd_data_bits_0_6; // @[Load.scala 97:29:@4945.4]
  assign io_inp_rd_data_bits_0_7 = tensorLoad_0_io_tensor_rd_data_bits_0_7; // @[Load.scala 97:29:@4946.4]
  assign io_inp_rd_data_bits_0_8 = tensorLoad_0_io_tensor_rd_data_bits_0_8; // @[Load.scala 97:29:@4947.4]
  assign io_inp_rd_data_bits_0_9 = tensorLoad_0_io_tensor_rd_data_bits_0_9; // @[Load.scala 97:29:@4948.4]
  assign io_inp_rd_data_bits_0_10 = tensorLoad_0_io_tensor_rd_data_bits_0_10; // @[Load.scala 97:29:@4949.4]
  assign io_inp_rd_data_bits_0_11 = tensorLoad_0_io_tensor_rd_data_bits_0_11; // @[Load.scala 97:29:@4950.4]
  assign io_inp_rd_data_bits_0_12 = tensorLoad_0_io_tensor_rd_data_bits_0_12; // @[Load.scala 97:29:@4951.4]
  assign io_inp_rd_data_bits_0_13 = tensorLoad_0_io_tensor_rd_data_bits_0_13; // @[Load.scala 97:29:@4952.4]
  assign io_inp_rd_data_bits_0_14 = tensorLoad_0_io_tensor_rd_data_bits_0_14; // @[Load.scala 97:29:@4953.4]
  assign io_inp_rd_data_bits_0_15 = tensorLoad_0_io_tensor_rd_data_bits_0_15; // @[Load.scala 97:29:@4954.4]
  assign io_wgt_rd_data_valid = tensorLoad_1_io_tensor_rd_data_valid; // @[Load.scala 97:29:@5485.4]
  assign io_wgt_rd_data_bits_0_0 = tensorLoad_1_io_tensor_rd_data_bits_0_0; // @[Load.scala 97:29:@5229.4]
  assign io_wgt_rd_data_bits_0_1 = tensorLoad_1_io_tensor_rd_data_bits_0_1; // @[Load.scala 97:29:@5230.4]
  assign io_wgt_rd_data_bits_0_2 = tensorLoad_1_io_tensor_rd_data_bits_0_2; // @[Load.scala 97:29:@5231.4]
  assign io_wgt_rd_data_bits_0_3 = tensorLoad_1_io_tensor_rd_data_bits_0_3; // @[Load.scala 97:29:@5232.4]
  assign io_wgt_rd_data_bits_0_4 = tensorLoad_1_io_tensor_rd_data_bits_0_4; // @[Load.scala 97:29:@5233.4]
  assign io_wgt_rd_data_bits_0_5 = tensorLoad_1_io_tensor_rd_data_bits_0_5; // @[Load.scala 97:29:@5234.4]
  assign io_wgt_rd_data_bits_0_6 = tensorLoad_1_io_tensor_rd_data_bits_0_6; // @[Load.scala 97:29:@5235.4]
  assign io_wgt_rd_data_bits_0_7 = tensorLoad_1_io_tensor_rd_data_bits_0_7; // @[Load.scala 97:29:@5236.4]
  assign io_wgt_rd_data_bits_0_8 = tensorLoad_1_io_tensor_rd_data_bits_0_8; // @[Load.scala 97:29:@5237.4]
  assign io_wgt_rd_data_bits_0_9 = tensorLoad_1_io_tensor_rd_data_bits_0_9; // @[Load.scala 97:29:@5238.4]
  assign io_wgt_rd_data_bits_0_10 = tensorLoad_1_io_tensor_rd_data_bits_0_10; // @[Load.scala 97:29:@5239.4]
  assign io_wgt_rd_data_bits_0_11 = tensorLoad_1_io_tensor_rd_data_bits_0_11; // @[Load.scala 97:29:@5240.4]
  assign io_wgt_rd_data_bits_0_12 = tensorLoad_1_io_tensor_rd_data_bits_0_12; // @[Load.scala 97:29:@5241.4]
  assign io_wgt_rd_data_bits_0_13 = tensorLoad_1_io_tensor_rd_data_bits_0_13; // @[Load.scala 97:29:@5242.4]
  assign io_wgt_rd_data_bits_0_14 = tensorLoad_1_io_tensor_rd_data_bits_0_14; // @[Load.scala 97:29:@5243.4]
  assign io_wgt_rd_data_bits_0_15 = tensorLoad_1_io_tensor_rd_data_bits_0_15; // @[Load.scala 97:29:@5244.4]
  assign io_wgt_rd_data_bits_1_0 = tensorLoad_1_io_tensor_rd_data_bits_1_0; // @[Load.scala 97:29:@5245.4]
  assign io_wgt_rd_data_bits_1_1 = tensorLoad_1_io_tensor_rd_data_bits_1_1; // @[Load.scala 97:29:@5246.4]
  assign io_wgt_rd_data_bits_1_2 = tensorLoad_1_io_tensor_rd_data_bits_1_2; // @[Load.scala 97:29:@5247.4]
  assign io_wgt_rd_data_bits_1_3 = tensorLoad_1_io_tensor_rd_data_bits_1_3; // @[Load.scala 97:29:@5248.4]
  assign io_wgt_rd_data_bits_1_4 = tensorLoad_1_io_tensor_rd_data_bits_1_4; // @[Load.scala 97:29:@5249.4]
  assign io_wgt_rd_data_bits_1_5 = tensorLoad_1_io_tensor_rd_data_bits_1_5; // @[Load.scala 97:29:@5250.4]
  assign io_wgt_rd_data_bits_1_6 = tensorLoad_1_io_tensor_rd_data_bits_1_6; // @[Load.scala 97:29:@5251.4]
  assign io_wgt_rd_data_bits_1_7 = tensorLoad_1_io_tensor_rd_data_bits_1_7; // @[Load.scala 97:29:@5252.4]
  assign io_wgt_rd_data_bits_1_8 = tensorLoad_1_io_tensor_rd_data_bits_1_8; // @[Load.scala 97:29:@5253.4]
  assign io_wgt_rd_data_bits_1_9 = tensorLoad_1_io_tensor_rd_data_bits_1_9; // @[Load.scala 97:29:@5254.4]
  assign io_wgt_rd_data_bits_1_10 = tensorLoad_1_io_tensor_rd_data_bits_1_10; // @[Load.scala 97:29:@5255.4]
  assign io_wgt_rd_data_bits_1_11 = tensorLoad_1_io_tensor_rd_data_bits_1_11; // @[Load.scala 97:29:@5256.4]
  assign io_wgt_rd_data_bits_1_12 = tensorLoad_1_io_tensor_rd_data_bits_1_12; // @[Load.scala 97:29:@5257.4]
  assign io_wgt_rd_data_bits_1_13 = tensorLoad_1_io_tensor_rd_data_bits_1_13; // @[Load.scala 97:29:@5258.4]
  assign io_wgt_rd_data_bits_1_14 = tensorLoad_1_io_tensor_rd_data_bits_1_14; // @[Load.scala 97:29:@5259.4]
  assign io_wgt_rd_data_bits_1_15 = tensorLoad_1_io_tensor_rd_data_bits_1_15; // @[Load.scala 97:29:@5260.4]
  assign io_wgt_rd_data_bits_2_0 = tensorLoad_1_io_tensor_rd_data_bits_2_0; // @[Load.scala 97:29:@5261.4]
  assign io_wgt_rd_data_bits_2_1 = tensorLoad_1_io_tensor_rd_data_bits_2_1; // @[Load.scala 97:29:@5262.4]
  assign io_wgt_rd_data_bits_2_2 = tensorLoad_1_io_tensor_rd_data_bits_2_2; // @[Load.scala 97:29:@5263.4]
  assign io_wgt_rd_data_bits_2_3 = tensorLoad_1_io_tensor_rd_data_bits_2_3; // @[Load.scala 97:29:@5264.4]
  assign io_wgt_rd_data_bits_2_4 = tensorLoad_1_io_tensor_rd_data_bits_2_4; // @[Load.scala 97:29:@5265.4]
  assign io_wgt_rd_data_bits_2_5 = tensorLoad_1_io_tensor_rd_data_bits_2_5; // @[Load.scala 97:29:@5266.4]
  assign io_wgt_rd_data_bits_2_6 = tensorLoad_1_io_tensor_rd_data_bits_2_6; // @[Load.scala 97:29:@5267.4]
  assign io_wgt_rd_data_bits_2_7 = tensorLoad_1_io_tensor_rd_data_bits_2_7; // @[Load.scala 97:29:@5268.4]
  assign io_wgt_rd_data_bits_2_8 = tensorLoad_1_io_tensor_rd_data_bits_2_8; // @[Load.scala 97:29:@5269.4]
  assign io_wgt_rd_data_bits_2_9 = tensorLoad_1_io_tensor_rd_data_bits_2_9; // @[Load.scala 97:29:@5270.4]
  assign io_wgt_rd_data_bits_2_10 = tensorLoad_1_io_tensor_rd_data_bits_2_10; // @[Load.scala 97:29:@5271.4]
  assign io_wgt_rd_data_bits_2_11 = tensorLoad_1_io_tensor_rd_data_bits_2_11; // @[Load.scala 97:29:@5272.4]
  assign io_wgt_rd_data_bits_2_12 = tensorLoad_1_io_tensor_rd_data_bits_2_12; // @[Load.scala 97:29:@5273.4]
  assign io_wgt_rd_data_bits_2_13 = tensorLoad_1_io_tensor_rd_data_bits_2_13; // @[Load.scala 97:29:@5274.4]
  assign io_wgt_rd_data_bits_2_14 = tensorLoad_1_io_tensor_rd_data_bits_2_14; // @[Load.scala 97:29:@5275.4]
  assign io_wgt_rd_data_bits_2_15 = tensorLoad_1_io_tensor_rd_data_bits_2_15; // @[Load.scala 97:29:@5276.4]
  assign io_wgt_rd_data_bits_3_0 = tensorLoad_1_io_tensor_rd_data_bits_3_0; // @[Load.scala 97:29:@5277.4]
  assign io_wgt_rd_data_bits_3_1 = tensorLoad_1_io_tensor_rd_data_bits_3_1; // @[Load.scala 97:29:@5278.4]
  assign io_wgt_rd_data_bits_3_2 = tensorLoad_1_io_tensor_rd_data_bits_3_2; // @[Load.scala 97:29:@5279.4]
  assign io_wgt_rd_data_bits_3_3 = tensorLoad_1_io_tensor_rd_data_bits_3_3; // @[Load.scala 97:29:@5280.4]
  assign io_wgt_rd_data_bits_3_4 = tensorLoad_1_io_tensor_rd_data_bits_3_4; // @[Load.scala 97:29:@5281.4]
  assign io_wgt_rd_data_bits_3_5 = tensorLoad_1_io_tensor_rd_data_bits_3_5; // @[Load.scala 97:29:@5282.4]
  assign io_wgt_rd_data_bits_3_6 = tensorLoad_1_io_tensor_rd_data_bits_3_6; // @[Load.scala 97:29:@5283.4]
  assign io_wgt_rd_data_bits_3_7 = tensorLoad_1_io_tensor_rd_data_bits_3_7; // @[Load.scala 97:29:@5284.4]
  assign io_wgt_rd_data_bits_3_8 = tensorLoad_1_io_tensor_rd_data_bits_3_8; // @[Load.scala 97:29:@5285.4]
  assign io_wgt_rd_data_bits_3_9 = tensorLoad_1_io_tensor_rd_data_bits_3_9; // @[Load.scala 97:29:@5286.4]
  assign io_wgt_rd_data_bits_3_10 = tensorLoad_1_io_tensor_rd_data_bits_3_10; // @[Load.scala 97:29:@5287.4]
  assign io_wgt_rd_data_bits_3_11 = tensorLoad_1_io_tensor_rd_data_bits_3_11; // @[Load.scala 97:29:@5288.4]
  assign io_wgt_rd_data_bits_3_12 = tensorLoad_1_io_tensor_rd_data_bits_3_12; // @[Load.scala 97:29:@5289.4]
  assign io_wgt_rd_data_bits_3_13 = tensorLoad_1_io_tensor_rd_data_bits_3_13; // @[Load.scala 97:29:@5290.4]
  assign io_wgt_rd_data_bits_3_14 = tensorLoad_1_io_tensor_rd_data_bits_3_14; // @[Load.scala 97:29:@5291.4]
  assign io_wgt_rd_data_bits_3_15 = tensorLoad_1_io_tensor_rd_data_bits_3_15; // @[Load.scala 97:29:@5292.4]
  assign io_wgt_rd_data_bits_4_0 = tensorLoad_1_io_tensor_rd_data_bits_4_0; // @[Load.scala 97:29:@5293.4]
  assign io_wgt_rd_data_bits_4_1 = tensorLoad_1_io_tensor_rd_data_bits_4_1; // @[Load.scala 97:29:@5294.4]
  assign io_wgt_rd_data_bits_4_2 = tensorLoad_1_io_tensor_rd_data_bits_4_2; // @[Load.scala 97:29:@5295.4]
  assign io_wgt_rd_data_bits_4_3 = tensorLoad_1_io_tensor_rd_data_bits_4_3; // @[Load.scala 97:29:@5296.4]
  assign io_wgt_rd_data_bits_4_4 = tensorLoad_1_io_tensor_rd_data_bits_4_4; // @[Load.scala 97:29:@5297.4]
  assign io_wgt_rd_data_bits_4_5 = tensorLoad_1_io_tensor_rd_data_bits_4_5; // @[Load.scala 97:29:@5298.4]
  assign io_wgt_rd_data_bits_4_6 = tensorLoad_1_io_tensor_rd_data_bits_4_6; // @[Load.scala 97:29:@5299.4]
  assign io_wgt_rd_data_bits_4_7 = tensorLoad_1_io_tensor_rd_data_bits_4_7; // @[Load.scala 97:29:@5300.4]
  assign io_wgt_rd_data_bits_4_8 = tensorLoad_1_io_tensor_rd_data_bits_4_8; // @[Load.scala 97:29:@5301.4]
  assign io_wgt_rd_data_bits_4_9 = tensorLoad_1_io_tensor_rd_data_bits_4_9; // @[Load.scala 97:29:@5302.4]
  assign io_wgt_rd_data_bits_4_10 = tensorLoad_1_io_tensor_rd_data_bits_4_10; // @[Load.scala 97:29:@5303.4]
  assign io_wgt_rd_data_bits_4_11 = tensorLoad_1_io_tensor_rd_data_bits_4_11; // @[Load.scala 97:29:@5304.4]
  assign io_wgt_rd_data_bits_4_12 = tensorLoad_1_io_tensor_rd_data_bits_4_12; // @[Load.scala 97:29:@5305.4]
  assign io_wgt_rd_data_bits_4_13 = tensorLoad_1_io_tensor_rd_data_bits_4_13; // @[Load.scala 97:29:@5306.4]
  assign io_wgt_rd_data_bits_4_14 = tensorLoad_1_io_tensor_rd_data_bits_4_14; // @[Load.scala 97:29:@5307.4]
  assign io_wgt_rd_data_bits_4_15 = tensorLoad_1_io_tensor_rd_data_bits_4_15; // @[Load.scala 97:29:@5308.4]
  assign io_wgt_rd_data_bits_5_0 = tensorLoad_1_io_tensor_rd_data_bits_5_0; // @[Load.scala 97:29:@5309.4]
  assign io_wgt_rd_data_bits_5_1 = tensorLoad_1_io_tensor_rd_data_bits_5_1; // @[Load.scala 97:29:@5310.4]
  assign io_wgt_rd_data_bits_5_2 = tensorLoad_1_io_tensor_rd_data_bits_5_2; // @[Load.scala 97:29:@5311.4]
  assign io_wgt_rd_data_bits_5_3 = tensorLoad_1_io_tensor_rd_data_bits_5_3; // @[Load.scala 97:29:@5312.4]
  assign io_wgt_rd_data_bits_5_4 = tensorLoad_1_io_tensor_rd_data_bits_5_4; // @[Load.scala 97:29:@5313.4]
  assign io_wgt_rd_data_bits_5_5 = tensorLoad_1_io_tensor_rd_data_bits_5_5; // @[Load.scala 97:29:@5314.4]
  assign io_wgt_rd_data_bits_5_6 = tensorLoad_1_io_tensor_rd_data_bits_5_6; // @[Load.scala 97:29:@5315.4]
  assign io_wgt_rd_data_bits_5_7 = tensorLoad_1_io_tensor_rd_data_bits_5_7; // @[Load.scala 97:29:@5316.4]
  assign io_wgt_rd_data_bits_5_8 = tensorLoad_1_io_tensor_rd_data_bits_5_8; // @[Load.scala 97:29:@5317.4]
  assign io_wgt_rd_data_bits_5_9 = tensorLoad_1_io_tensor_rd_data_bits_5_9; // @[Load.scala 97:29:@5318.4]
  assign io_wgt_rd_data_bits_5_10 = tensorLoad_1_io_tensor_rd_data_bits_5_10; // @[Load.scala 97:29:@5319.4]
  assign io_wgt_rd_data_bits_5_11 = tensorLoad_1_io_tensor_rd_data_bits_5_11; // @[Load.scala 97:29:@5320.4]
  assign io_wgt_rd_data_bits_5_12 = tensorLoad_1_io_tensor_rd_data_bits_5_12; // @[Load.scala 97:29:@5321.4]
  assign io_wgt_rd_data_bits_5_13 = tensorLoad_1_io_tensor_rd_data_bits_5_13; // @[Load.scala 97:29:@5322.4]
  assign io_wgt_rd_data_bits_5_14 = tensorLoad_1_io_tensor_rd_data_bits_5_14; // @[Load.scala 97:29:@5323.4]
  assign io_wgt_rd_data_bits_5_15 = tensorLoad_1_io_tensor_rd_data_bits_5_15; // @[Load.scala 97:29:@5324.4]
  assign io_wgt_rd_data_bits_6_0 = tensorLoad_1_io_tensor_rd_data_bits_6_0; // @[Load.scala 97:29:@5325.4]
  assign io_wgt_rd_data_bits_6_1 = tensorLoad_1_io_tensor_rd_data_bits_6_1; // @[Load.scala 97:29:@5326.4]
  assign io_wgt_rd_data_bits_6_2 = tensorLoad_1_io_tensor_rd_data_bits_6_2; // @[Load.scala 97:29:@5327.4]
  assign io_wgt_rd_data_bits_6_3 = tensorLoad_1_io_tensor_rd_data_bits_6_3; // @[Load.scala 97:29:@5328.4]
  assign io_wgt_rd_data_bits_6_4 = tensorLoad_1_io_tensor_rd_data_bits_6_4; // @[Load.scala 97:29:@5329.4]
  assign io_wgt_rd_data_bits_6_5 = tensorLoad_1_io_tensor_rd_data_bits_6_5; // @[Load.scala 97:29:@5330.4]
  assign io_wgt_rd_data_bits_6_6 = tensorLoad_1_io_tensor_rd_data_bits_6_6; // @[Load.scala 97:29:@5331.4]
  assign io_wgt_rd_data_bits_6_7 = tensorLoad_1_io_tensor_rd_data_bits_6_7; // @[Load.scala 97:29:@5332.4]
  assign io_wgt_rd_data_bits_6_8 = tensorLoad_1_io_tensor_rd_data_bits_6_8; // @[Load.scala 97:29:@5333.4]
  assign io_wgt_rd_data_bits_6_9 = tensorLoad_1_io_tensor_rd_data_bits_6_9; // @[Load.scala 97:29:@5334.4]
  assign io_wgt_rd_data_bits_6_10 = tensorLoad_1_io_tensor_rd_data_bits_6_10; // @[Load.scala 97:29:@5335.4]
  assign io_wgt_rd_data_bits_6_11 = tensorLoad_1_io_tensor_rd_data_bits_6_11; // @[Load.scala 97:29:@5336.4]
  assign io_wgt_rd_data_bits_6_12 = tensorLoad_1_io_tensor_rd_data_bits_6_12; // @[Load.scala 97:29:@5337.4]
  assign io_wgt_rd_data_bits_6_13 = tensorLoad_1_io_tensor_rd_data_bits_6_13; // @[Load.scala 97:29:@5338.4]
  assign io_wgt_rd_data_bits_6_14 = tensorLoad_1_io_tensor_rd_data_bits_6_14; // @[Load.scala 97:29:@5339.4]
  assign io_wgt_rd_data_bits_6_15 = tensorLoad_1_io_tensor_rd_data_bits_6_15; // @[Load.scala 97:29:@5340.4]
  assign io_wgt_rd_data_bits_7_0 = tensorLoad_1_io_tensor_rd_data_bits_7_0; // @[Load.scala 97:29:@5341.4]
  assign io_wgt_rd_data_bits_7_1 = tensorLoad_1_io_tensor_rd_data_bits_7_1; // @[Load.scala 97:29:@5342.4]
  assign io_wgt_rd_data_bits_7_2 = tensorLoad_1_io_tensor_rd_data_bits_7_2; // @[Load.scala 97:29:@5343.4]
  assign io_wgt_rd_data_bits_7_3 = tensorLoad_1_io_tensor_rd_data_bits_7_3; // @[Load.scala 97:29:@5344.4]
  assign io_wgt_rd_data_bits_7_4 = tensorLoad_1_io_tensor_rd_data_bits_7_4; // @[Load.scala 97:29:@5345.4]
  assign io_wgt_rd_data_bits_7_5 = tensorLoad_1_io_tensor_rd_data_bits_7_5; // @[Load.scala 97:29:@5346.4]
  assign io_wgt_rd_data_bits_7_6 = tensorLoad_1_io_tensor_rd_data_bits_7_6; // @[Load.scala 97:29:@5347.4]
  assign io_wgt_rd_data_bits_7_7 = tensorLoad_1_io_tensor_rd_data_bits_7_7; // @[Load.scala 97:29:@5348.4]
  assign io_wgt_rd_data_bits_7_8 = tensorLoad_1_io_tensor_rd_data_bits_7_8; // @[Load.scala 97:29:@5349.4]
  assign io_wgt_rd_data_bits_7_9 = tensorLoad_1_io_tensor_rd_data_bits_7_9; // @[Load.scala 97:29:@5350.4]
  assign io_wgt_rd_data_bits_7_10 = tensorLoad_1_io_tensor_rd_data_bits_7_10; // @[Load.scala 97:29:@5351.4]
  assign io_wgt_rd_data_bits_7_11 = tensorLoad_1_io_tensor_rd_data_bits_7_11; // @[Load.scala 97:29:@5352.4]
  assign io_wgt_rd_data_bits_7_12 = tensorLoad_1_io_tensor_rd_data_bits_7_12; // @[Load.scala 97:29:@5353.4]
  assign io_wgt_rd_data_bits_7_13 = tensorLoad_1_io_tensor_rd_data_bits_7_13; // @[Load.scala 97:29:@5354.4]
  assign io_wgt_rd_data_bits_7_14 = tensorLoad_1_io_tensor_rd_data_bits_7_14; // @[Load.scala 97:29:@5355.4]
  assign io_wgt_rd_data_bits_7_15 = tensorLoad_1_io_tensor_rd_data_bits_7_15; // @[Load.scala 97:29:@5356.4]
  assign io_wgt_rd_data_bits_8_0 = tensorLoad_1_io_tensor_rd_data_bits_8_0; // @[Load.scala 97:29:@5357.4]
  assign io_wgt_rd_data_bits_8_1 = tensorLoad_1_io_tensor_rd_data_bits_8_1; // @[Load.scala 97:29:@5358.4]
  assign io_wgt_rd_data_bits_8_2 = tensorLoad_1_io_tensor_rd_data_bits_8_2; // @[Load.scala 97:29:@5359.4]
  assign io_wgt_rd_data_bits_8_3 = tensorLoad_1_io_tensor_rd_data_bits_8_3; // @[Load.scala 97:29:@5360.4]
  assign io_wgt_rd_data_bits_8_4 = tensorLoad_1_io_tensor_rd_data_bits_8_4; // @[Load.scala 97:29:@5361.4]
  assign io_wgt_rd_data_bits_8_5 = tensorLoad_1_io_tensor_rd_data_bits_8_5; // @[Load.scala 97:29:@5362.4]
  assign io_wgt_rd_data_bits_8_6 = tensorLoad_1_io_tensor_rd_data_bits_8_6; // @[Load.scala 97:29:@5363.4]
  assign io_wgt_rd_data_bits_8_7 = tensorLoad_1_io_tensor_rd_data_bits_8_7; // @[Load.scala 97:29:@5364.4]
  assign io_wgt_rd_data_bits_8_8 = tensorLoad_1_io_tensor_rd_data_bits_8_8; // @[Load.scala 97:29:@5365.4]
  assign io_wgt_rd_data_bits_8_9 = tensorLoad_1_io_tensor_rd_data_bits_8_9; // @[Load.scala 97:29:@5366.4]
  assign io_wgt_rd_data_bits_8_10 = tensorLoad_1_io_tensor_rd_data_bits_8_10; // @[Load.scala 97:29:@5367.4]
  assign io_wgt_rd_data_bits_8_11 = tensorLoad_1_io_tensor_rd_data_bits_8_11; // @[Load.scala 97:29:@5368.4]
  assign io_wgt_rd_data_bits_8_12 = tensorLoad_1_io_tensor_rd_data_bits_8_12; // @[Load.scala 97:29:@5369.4]
  assign io_wgt_rd_data_bits_8_13 = tensorLoad_1_io_tensor_rd_data_bits_8_13; // @[Load.scala 97:29:@5370.4]
  assign io_wgt_rd_data_bits_8_14 = tensorLoad_1_io_tensor_rd_data_bits_8_14; // @[Load.scala 97:29:@5371.4]
  assign io_wgt_rd_data_bits_8_15 = tensorLoad_1_io_tensor_rd_data_bits_8_15; // @[Load.scala 97:29:@5372.4]
  assign io_wgt_rd_data_bits_9_0 = tensorLoad_1_io_tensor_rd_data_bits_9_0; // @[Load.scala 97:29:@5373.4]
  assign io_wgt_rd_data_bits_9_1 = tensorLoad_1_io_tensor_rd_data_bits_9_1; // @[Load.scala 97:29:@5374.4]
  assign io_wgt_rd_data_bits_9_2 = tensorLoad_1_io_tensor_rd_data_bits_9_2; // @[Load.scala 97:29:@5375.4]
  assign io_wgt_rd_data_bits_9_3 = tensorLoad_1_io_tensor_rd_data_bits_9_3; // @[Load.scala 97:29:@5376.4]
  assign io_wgt_rd_data_bits_9_4 = tensorLoad_1_io_tensor_rd_data_bits_9_4; // @[Load.scala 97:29:@5377.4]
  assign io_wgt_rd_data_bits_9_5 = tensorLoad_1_io_tensor_rd_data_bits_9_5; // @[Load.scala 97:29:@5378.4]
  assign io_wgt_rd_data_bits_9_6 = tensorLoad_1_io_tensor_rd_data_bits_9_6; // @[Load.scala 97:29:@5379.4]
  assign io_wgt_rd_data_bits_9_7 = tensorLoad_1_io_tensor_rd_data_bits_9_7; // @[Load.scala 97:29:@5380.4]
  assign io_wgt_rd_data_bits_9_8 = tensorLoad_1_io_tensor_rd_data_bits_9_8; // @[Load.scala 97:29:@5381.4]
  assign io_wgt_rd_data_bits_9_9 = tensorLoad_1_io_tensor_rd_data_bits_9_9; // @[Load.scala 97:29:@5382.4]
  assign io_wgt_rd_data_bits_9_10 = tensorLoad_1_io_tensor_rd_data_bits_9_10; // @[Load.scala 97:29:@5383.4]
  assign io_wgt_rd_data_bits_9_11 = tensorLoad_1_io_tensor_rd_data_bits_9_11; // @[Load.scala 97:29:@5384.4]
  assign io_wgt_rd_data_bits_9_12 = tensorLoad_1_io_tensor_rd_data_bits_9_12; // @[Load.scala 97:29:@5385.4]
  assign io_wgt_rd_data_bits_9_13 = tensorLoad_1_io_tensor_rd_data_bits_9_13; // @[Load.scala 97:29:@5386.4]
  assign io_wgt_rd_data_bits_9_14 = tensorLoad_1_io_tensor_rd_data_bits_9_14; // @[Load.scala 97:29:@5387.4]
  assign io_wgt_rd_data_bits_9_15 = tensorLoad_1_io_tensor_rd_data_bits_9_15; // @[Load.scala 97:29:@5388.4]
  assign io_wgt_rd_data_bits_10_0 = tensorLoad_1_io_tensor_rd_data_bits_10_0; // @[Load.scala 97:29:@5389.4]
  assign io_wgt_rd_data_bits_10_1 = tensorLoad_1_io_tensor_rd_data_bits_10_1; // @[Load.scala 97:29:@5390.4]
  assign io_wgt_rd_data_bits_10_2 = tensorLoad_1_io_tensor_rd_data_bits_10_2; // @[Load.scala 97:29:@5391.4]
  assign io_wgt_rd_data_bits_10_3 = tensorLoad_1_io_tensor_rd_data_bits_10_3; // @[Load.scala 97:29:@5392.4]
  assign io_wgt_rd_data_bits_10_4 = tensorLoad_1_io_tensor_rd_data_bits_10_4; // @[Load.scala 97:29:@5393.4]
  assign io_wgt_rd_data_bits_10_5 = tensorLoad_1_io_tensor_rd_data_bits_10_5; // @[Load.scala 97:29:@5394.4]
  assign io_wgt_rd_data_bits_10_6 = tensorLoad_1_io_tensor_rd_data_bits_10_6; // @[Load.scala 97:29:@5395.4]
  assign io_wgt_rd_data_bits_10_7 = tensorLoad_1_io_tensor_rd_data_bits_10_7; // @[Load.scala 97:29:@5396.4]
  assign io_wgt_rd_data_bits_10_8 = tensorLoad_1_io_tensor_rd_data_bits_10_8; // @[Load.scala 97:29:@5397.4]
  assign io_wgt_rd_data_bits_10_9 = tensorLoad_1_io_tensor_rd_data_bits_10_9; // @[Load.scala 97:29:@5398.4]
  assign io_wgt_rd_data_bits_10_10 = tensorLoad_1_io_tensor_rd_data_bits_10_10; // @[Load.scala 97:29:@5399.4]
  assign io_wgt_rd_data_bits_10_11 = tensorLoad_1_io_tensor_rd_data_bits_10_11; // @[Load.scala 97:29:@5400.4]
  assign io_wgt_rd_data_bits_10_12 = tensorLoad_1_io_tensor_rd_data_bits_10_12; // @[Load.scala 97:29:@5401.4]
  assign io_wgt_rd_data_bits_10_13 = tensorLoad_1_io_tensor_rd_data_bits_10_13; // @[Load.scala 97:29:@5402.4]
  assign io_wgt_rd_data_bits_10_14 = tensorLoad_1_io_tensor_rd_data_bits_10_14; // @[Load.scala 97:29:@5403.4]
  assign io_wgt_rd_data_bits_10_15 = tensorLoad_1_io_tensor_rd_data_bits_10_15; // @[Load.scala 97:29:@5404.4]
  assign io_wgt_rd_data_bits_11_0 = tensorLoad_1_io_tensor_rd_data_bits_11_0; // @[Load.scala 97:29:@5405.4]
  assign io_wgt_rd_data_bits_11_1 = tensorLoad_1_io_tensor_rd_data_bits_11_1; // @[Load.scala 97:29:@5406.4]
  assign io_wgt_rd_data_bits_11_2 = tensorLoad_1_io_tensor_rd_data_bits_11_2; // @[Load.scala 97:29:@5407.4]
  assign io_wgt_rd_data_bits_11_3 = tensorLoad_1_io_tensor_rd_data_bits_11_3; // @[Load.scala 97:29:@5408.4]
  assign io_wgt_rd_data_bits_11_4 = tensorLoad_1_io_tensor_rd_data_bits_11_4; // @[Load.scala 97:29:@5409.4]
  assign io_wgt_rd_data_bits_11_5 = tensorLoad_1_io_tensor_rd_data_bits_11_5; // @[Load.scala 97:29:@5410.4]
  assign io_wgt_rd_data_bits_11_6 = tensorLoad_1_io_tensor_rd_data_bits_11_6; // @[Load.scala 97:29:@5411.4]
  assign io_wgt_rd_data_bits_11_7 = tensorLoad_1_io_tensor_rd_data_bits_11_7; // @[Load.scala 97:29:@5412.4]
  assign io_wgt_rd_data_bits_11_8 = tensorLoad_1_io_tensor_rd_data_bits_11_8; // @[Load.scala 97:29:@5413.4]
  assign io_wgt_rd_data_bits_11_9 = tensorLoad_1_io_tensor_rd_data_bits_11_9; // @[Load.scala 97:29:@5414.4]
  assign io_wgt_rd_data_bits_11_10 = tensorLoad_1_io_tensor_rd_data_bits_11_10; // @[Load.scala 97:29:@5415.4]
  assign io_wgt_rd_data_bits_11_11 = tensorLoad_1_io_tensor_rd_data_bits_11_11; // @[Load.scala 97:29:@5416.4]
  assign io_wgt_rd_data_bits_11_12 = tensorLoad_1_io_tensor_rd_data_bits_11_12; // @[Load.scala 97:29:@5417.4]
  assign io_wgt_rd_data_bits_11_13 = tensorLoad_1_io_tensor_rd_data_bits_11_13; // @[Load.scala 97:29:@5418.4]
  assign io_wgt_rd_data_bits_11_14 = tensorLoad_1_io_tensor_rd_data_bits_11_14; // @[Load.scala 97:29:@5419.4]
  assign io_wgt_rd_data_bits_11_15 = tensorLoad_1_io_tensor_rd_data_bits_11_15; // @[Load.scala 97:29:@5420.4]
  assign io_wgt_rd_data_bits_12_0 = tensorLoad_1_io_tensor_rd_data_bits_12_0; // @[Load.scala 97:29:@5421.4]
  assign io_wgt_rd_data_bits_12_1 = tensorLoad_1_io_tensor_rd_data_bits_12_1; // @[Load.scala 97:29:@5422.4]
  assign io_wgt_rd_data_bits_12_2 = tensorLoad_1_io_tensor_rd_data_bits_12_2; // @[Load.scala 97:29:@5423.4]
  assign io_wgt_rd_data_bits_12_3 = tensorLoad_1_io_tensor_rd_data_bits_12_3; // @[Load.scala 97:29:@5424.4]
  assign io_wgt_rd_data_bits_12_4 = tensorLoad_1_io_tensor_rd_data_bits_12_4; // @[Load.scala 97:29:@5425.4]
  assign io_wgt_rd_data_bits_12_5 = tensorLoad_1_io_tensor_rd_data_bits_12_5; // @[Load.scala 97:29:@5426.4]
  assign io_wgt_rd_data_bits_12_6 = tensorLoad_1_io_tensor_rd_data_bits_12_6; // @[Load.scala 97:29:@5427.4]
  assign io_wgt_rd_data_bits_12_7 = tensorLoad_1_io_tensor_rd_data_bits_12_7; // @[Load.scala 97:29:@5428.4]
  assign io_wgt_rd_data_bits_12_8 = tensorLoad_1_io_tensor_rd_data_bits_12_8; // @[Load.scala 97:29:@5429.4]
  assign io_wgt_rd_data_bits_12_9 = tensorLoad_1_io_tensor_rd_data_bits_12_9; // @[Load.scala 97:29:@5430.4]
  assign io_wgt_rd_data_bits_12_10 = tensorLoad_1_io_tensor_rd_data_bits_12_10; // @[Load.scala 97:29:@5431.4]
  assign io_wgt_rd_data_bits_12_11 = tensorLoad_1_io_tensor_rd_data_bits_12_11; // @[Load.scala 97:29:@5432.4]
  assign io_wgt_rd_data_bits_12_12 = tensorLoad_1_io_tensor_rd_data_bits_12_12; // @[Load.scala 97:29:@5433.4]
  assign io_wgt_rd_data_bits_12_13 = tensorLoad_1_io_tensor_rd_data_bits_12_13; // @[Load.scala 97:29:@5434.4]
  assign io_wgt_rd_data_bits_12_14 = tensorLoad_1_io_tensor_rd_data_bits_12_14; // @[Load.scala 97:29:@5435.4]
  assign io_wgt_rd_data_bits_12_15 = tensorLoad_1_io_tensor_rd_data_bits_12_15; // @[Load.scala 97:29:@5436.4]
  assign io_wgt_rd_data_bits_13_0 = tensorLoad_1_io_tensor_rd_data_bits_13_0; // @[Load.scala 97:29:@5437.4]
  assign io_wgt_rd_data_bits_13_1 = tensorLoad_1_io_tensor_rd_data_bits_13_1; // @[Load.scala 97:29:@5438.4]
  assign io_wgt_rd_data_bits_13_2 = tensorLoad_1_io_tensor_rd_data_bits_13_2; // @[Load.scala 97:29:@5439.4]
  assign io_wgt_rd_data_bits_13_3 = tensorLoad_1_io_tensor_rd_data_bits_13_3; // @[Load.scala 97:29:@5440.4]
  assign io_wgt_rd_data_bits_13_4 = tensorLoad_1_io_tensor_rd_data_bits_13_4; // @[Load.scala 97:29:@5441.4]
  assign io_wgt_rd_data_bits_13_5 = tensorLoad_1_io_tensor_rd_data_bits_13_5; // @[Load.scala 97:29:@5442.4]
  assign io_wgt_rd_data_bits_13_6 = tensorLoad_1_io_tensor_rd_data_bits_13_6; // @[Load.scala 97:29:@5443.4]
  assign io_wgt_rd_data_bits_13_7 = tensorLoad_1_io_tensor_rd_data_bits_13_7; // @[Load.scala 97:29:@5444.4]
  assign io_wgt_rd_data_bits_13_8 = tensorLoad_1_io_tensor_rd_data_bits_13_8; // @[Load.scala 97:29:@5445.4]
  assign io_wgt_rd_data_bits_13_9 = tensorLoad_1_io_tensor_rd_data_bits_13_9; // @[Load.scala 97:29:@5446.4]
  assign io_wgt_rd_data_bits_13_10 = tensorLoad_1_io_tensor_rd_data_bits_13_10; // @[Load.scala 97:29:@5447.4]
  assign io_wgt_rd_data_bits_13_11 = tensorLoad_1_io_tensor_rd_data_bits_13_11; // @[Load.scala 97:29:@5448.4]
  assign io_wgt_rd_data_bits_13_12 = tensorLoad_1_io_tensor_rd_data_bits_13_12; // @[Load.scala 97:29:@5449.4]
  assign io_wgt_rd_data_bits_13_13 = tensorLoad_1_io_tensor_rd_data_bits_13_13; // @[Load.scala 97:29:@5450.4]
  assign io_wgt_rd_data_bits_13_14 = tensorLoad_1_io_tensor_rd_data_bits_13_14; // @[Load.scala 97:29:@5451.4]
  assign io_wgt_rd_data_bits_13_15 = tensorLoad_1_io_tensor_rd_data_bits_13_15; // @[Load.scala 97:29:@5452.4]
  assign io_wgt_rd_data_bits_14_0 = tensorLoad_1_io_tensor_rd_data_bits_14_0; // @[Load.scala 97:29:@5453.4]
  assign io_wgt_rd_data_bits_14_1 = tensorLoad_1_io_tensor_rd_data_bits_14_1; // @[Load.scala 97:29:@5454.4]
  assign io_wgt_rd_data_bits_14_2 = tensorLoad_1_io_tensor_rd_data_bits_14_2; // @[Load.scala 97:29:@5455.4]
  assign io_wgt_rd_data_bits_14_3 = tensorLoad_1_io_tensor_rd_data_bits_14_3; // @[Load.scala 97:29:@5456.4]
  assign io_wgt_rd_data_bits_14_4 = tensorLoad_1_io_tensor_rd_data_bits_14_4; // @[Load.scala 97:29:@5457.4]
  assign io_wgt_rd_data_bits_14_5 = tensorLoad_1_io_tensor_rd_data_bits_14_5; // @[Load.scala 97:29:@5458.4]
  assign io_wgt_rd_data_bits_14_6 = tensorLoad_1_io_tensor_rd_data_bits_14_6; // @[Load.scala 97:29:@5459.4]
  assign io_wgt_rd_data_bits_14_7 = tensorLoad_1_io_tensor_rd_data_bits_14_7; // @[Load.scala 97:29:@5460.4]
  assign io_wgt_rd_data_bits_14_8 = tensorLoad_1_io_tensor_rd_data_bits_14_8; // @[Load.scala 97:29:@5461.4]
  assign io_wgt_rd_data_bits_14_9 = tensorLoad_1_io_tensor_rd_data_bits_14_9; // @[Load.scala 97:29:@5462.4]
  assign io_wgt_rd_data_bits_14_10 = tensorLoad_1_io_tensor_rd_data_bits_14_10; // @[Load.scala 97:29:@5463.4]
  assign io_wgt_rd_data_bits_14_11 = tensorLoad_1_io_tensor_rd_data_bits_14_11; // @[Load.scala 97:29:@5464.4]
  assign io_wgt_rd_data_bits_14_12 = tensorLoad_1_io_tensor_rd_data_bits_14_12; // @[Load.scala 97:29:@5465.4]
  assign io_wgt_rd_data_bits_14_13 = tensorLoad_1_io_tensor_rd_data_bits_14_13; // @[Load.scala 97:29:@5466.4]
  assign io_wgt_rd_data_bits_14_14 = tensorLoad_1_io_tensor_rd_data_bits_14_14; // @[Load.scala 97:29:@5467.4]
  assign io_wgt_rd_data_bits_14_15 = tensorLoad_1_io_tensor_rd_data_bits_14_15; // @[Load.scala 97:29:@5468.4]
  assign io_wgt_rd_data_bits_15_0 = tensorLoad_1_io_tensor_rd_data_bits_15_0; // @[Load.scala 97:29:@5469.4]
  assign io_wgt_rd_data_bits_15_1 = tensorLoad_1_io_tensor_rd_data_bits_15_1; // @[Load.scala 97:29:@5470.4]
  assign io_wgt_rd_data_bits_15_2 = tensorLoad_1_io_tensor_rd_data_bits_15_2; // @[Load.scala 97:29:@5471.4]
  assign io_wgt_rd_data_bits_15_3 = tensorLoad_1_io_tensor_rd_data_bits_15_3; // @[Load.scala 97:29:@5472.4]
  assign io_wgt_rd_data_bits_15_4 = tensorLoad_1_io_tensor_rd_data_bits_15_4; // @[Load.scala 97:29:@5473.4]
  assign io_wgt_rd_data_bits_15_5 = tensorLoad_1_io_tensor_rd_data_bits_15_5; // @[Load.scala 97:29:@5474.4]
  assign io_wgt_rd_data_bits_15_6 = tensorLoad_1_io_tensor_rd_data_bits_15_6; // @[Load.scala 97:29:@5475.4]
  assign io_wgt_rd_data_bits_15_7 = tensorLoad_1_io_tensor_rd_data_bits_15_7; // @[Load.scala 97:29:@5476.4]
  assign io_wgt_rd_data_bits_15_8 = tensorLoad_1_io_tensor_rd_data_bits_15_8; // @[Load.scala 97:29:@5477.4]
  assign io_wgt_rd_data_bits_15_9 = tensorLoad_1_io_tensor_rd_data_bits_15_9; // @[Load.scala 97:29:@5478.4]
  assign io_wgt_rd_data_bits_15_10 = tensorLoad_1_io_tensor_rd_data_bits_15_10; // @[Load.scala 97:29:@5479.4]
  assign io_wgt_rd_data_bits_15_11 = tensorLoad_1_io_tensor_rd_data_bits_15_11; // @[Load.scala 97:29:@5480.4]
  assign io_wgt_rd_data_bits_15_12 = tensorLoad_1_io_tensor_rd_data_bits_15_12; // @[Load.scala 97:29:@5481.4]
  assign io_wgt_rd_data_bits_15_13 = tensorLoad_1_io_tensor_rd_data_bits_15_13; // @[Load.scala 97:29:@5482.4]
  assign io_wgt_rd_data_bits_15_14 = tensorLoad_1_io_tensor_rd_data_bits_15_14; // @[Load.scala 97:29:@5483.4]
  assign io_wgt_rd_data_bits_15_15 = tensorLoad_1_io_tensor_rd_data_bits_15_15; // @[Load.scala 97:29:@5484.4]
  assign s_clock = clock; // @[:@4864.4]
  assign s_reset = reset; // @[:@4865.4]
  assign s_io_spost = io_i_post; // @[Load.scala 102:14:@5495.4]
  assign s_io_swait = dec_io_pop_next & _T_5009; // @[Load.scala 103:14:@5499.4]
  assign inst_q_clock = clock; // @[:@4867.4]
  assign inst_q_reset = reset; // @[:@4868.4]
  assign inst_q_io_enq_valid = io_inst_valid; // @[Load.scala 85:17:@4908.4]
  assign inst_q_io_enq_bits = io_inst_bits; // @[Load.scala 85:17:@4907.4]
  assign inst_q_io_deq_ready = _T_5005 | _T_5006; // @[Load.scala 86:23:@4914.4]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Load.scala 53:15:@4872.4]
  assign tensorLoad_0_clock = clock; // @[:@4874.4]
  assign tensorLoad_0_reset = reset; // @[:@4875.4]
  assign tensorLoad_0_io_start = _T_5009 & dec_io_isInput; // @[Load.scala 94:28:@4918.4]
  assign tensorLoad_0_io_inst = inst_q_io_deq_bits; // @[Load.scala 95:27:@4919.4]
  assign tensorLoad_0_io_baddr = io_inp_baddr; // @[Load.scala 96:28:@4920.4]
  assign tensorLoad_0_io_vme_rd_cmd_ready = io_vme_rd_0_cmd_ready; // @[Load.scala 98:18:@4964.4]
  assign tensorLoad_0_io_vme_rd_data_valid = io_vme_rd_0_data_valid; // @[Load.scala 98:18:@4959.4]
  assign tensorLoad_0_io_vme_rd_data_bits = io_vme_rd_0_data_bits; // @[Load.scala 98:18:@4958.4]
  assign tensorLoad_0_io_tensor_rd_idx_valid = io_inp_rd_idx_valid; // @[Load.scala 97:29:@4957.4]
  assign tensorLoad_0_io_tensor_rd_idx_bits = io_inp_rd_idx_bits; // @[Load.scala 97:29:@4956.4]
  assign tensorLoad_1_clock = clock; // @[:@4877.4]
  assign tensorLoad_1_reset = reset; // @[:@4878.4]
  assign tensorLoad_1_io_start = _T_5009 & dec_io_isWeight; // @[Load.scala 94:28:@4968.4]
  assign tensorLoad_1_io_inst = inst_q_io_deq_bits; // @[Load.scala 95:27:@4969.4]
  assign tensorLoad_1_io_baddr = io_wgt_baddr; // @[Load.scala 96:28:@4970.4]
  assign tensorLoad_1_io_vme_rd_cmd_ready = io_vme_rd_1_cmd_ready; // @[Load.scala 98:18:@5494.4]
  assign tensorLoad_1_io_vme_rd_data_valid = io_vme_rd_1_data_valid; // @[Load.scala 98:18:@5489.4]
  assign tensorLoad_1_io_vme_rd_data_bits = io_vme_rd_1_data_bits; // @[Load.scala 98:18:@5488.4]
  assign tensorLoad_1_io_tensor_rd_idx_valid = io_wgt_rd_idx_valid; // @[Load.scala 97:29:@5487.4]
  assign tensorLoad_1_io_tensor_rd_idx_bits = io_wgt_rd_idx_bits; // @[Load.scala 97:29:@5486.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_5000) begin
        if (start) begin
          if (dec_io_isSync) begin
            state <= 2'h1;
          end else begin
            if (_T_5001) begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_5002) begin
          state <= 2'h0;
        end else begin
          if (_T_5003) begin
            if (done) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module LoadUop( // @[:@5563.2]
  input          clock, // @[:@5564.4]
  input          reset, // @[:@5565.4]
  input          io_start, // @[:@5566.4]
  output         io_done, // @[:@5566.4]
  input  [127:0] io_inst, // @[:@5566.4]
  input  [31:0]  io_baddr, // @[:@5566.4]
  input          io_vme_rd_cmd_ready, // @[:@5566.4]
  output         io_vme_rd_cmd_valid, // @[:@5566.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@5566.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@5566.4]
  output         io_vme_rd_data_ready, // @[:@5566.4]
  input          io_vme_rd_data_valid, // @[:@5566.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@5566.4]
  input          io_uop_idx_valid, // @[:@5566.4]
  input  [10:0]  io_uop_idx_bits, // @[:@5566.4]
  output         io_uop_data_valid, // @[:@5566.4]
  output [9:0]   io_uop_data_bits_u2, // @[:@5566.4]
  output [10:0]  io_uop_data_bits_u1, // @[:@5566.4]
  output [10:0]  io_uop_data_bits_u0 // @[:@5566.4]
);
  reg [31:0] mem_0 [0:1023]; // @[LoadUop.scala 163:24:@5800.4]
  reg [31:0] _RAND_0;
  wire [31:0] mem_0_memRead_data; // @[LoadUop.scala 163:24:@5800.4]
  wire [9:0] mem_0_memRead_addr; // @[LoadUop.scala 163:24:@5800.4]
  wire [31:0] mem_0__T_564_data; // @[LoadUop.scala 163:24:@5800.4]
  wire [9:0] mem_0__T_564_addr; // @[LoadUop.scala 163:24:@5800.4]
  wire  mem_0__T_564_mask; // @[LoadUop.scala 163:24:@5800.4]
  wire  mem_0__T_564_en; // @[LoadUop.scala 163:24:@5800.4]
  reg [31:0] mem_1 [0:1023]; // @[LoadUop.scala 163:24:@5800.4]
  reg [31:0] _RAND_1;
  wire [31:0] mem_1_memRead_data; // @[LoadUop.scala 163:24:@5800.4]
  wire [9:0] mem_1_memRead_addr; // @[LoadUop.scala 163:24:@5800.4]
  wire [31:0] mem_1__T_564_data; // @[LoadUop.scala 163:24:@5800.4]
  wire [9:0] mem_1__T_564_addr; // @[LoadUop.scala 163:24:@5800.4]
  wire  mem_1__T_564_mask; // @[LoadUop.scala 163:24:@5800.4]
  wire  mem_1__T_564_en; // @[LoadUop.scala 163:24:@5800.4]
  wire [15:0] dec_sram_offset; // @[LoadUop.scala 75:29:@5583.4]
  wire [31:0] dec_dram_offset; // @[LoadUop.scala 75:29:@5585.4]
  wire [15:0] dec_xsize; // @[LoadUop.scala 75:29:@5591.4]
  reg [31:0] raddr; // @[LoadUop.scala 76:18:@5603.4]
  reg [31:0] _RAND_2;
  reg [7:0] xcnt; // @[LoadUop.scala 77:17:@5604.4]
  reg [31:0] _RAND_3;
  reg [7:0] xlen; // @[LoadUop.scala 78:17:@5605.4]
  reg [31:0] _RAND_4;
  reg [15:0] xrem; // @[LoadUop.scala 79:17:@5606.4]
  reg [31:0] _RAND_5;
  wire [14:0] _T_67; // @[LoadUop.scala 80:26:@5607.4]
  wire  _T_68; // @[LoadUop.scala 80:58:@5608.4]
  wire [14:0] _GEN_89; // @[LoadUop.scala 80:47:@5609.4]
  wire [15:0] _T_69; // @[LoadUop.scala 80:47:@5609.4]
  wire [14:0] _T_70; // @[LoadUop.scala 80:47:@5610.4]
  wire [15:0] _GEN_6; // @[LoadUop.scala 80:81:@5611.4]
  wire [1:0] _T_72; // @[LoadUop.scala 80:81:@5611.4]
  wire [14:0] _GEN_90; // @[LoadUop.scala 80:62:@5612.4]
  wire [15:0] _T_73; // @[LoadUop.scala 80:62:@5612.4]
  wire [14:0] _T_74; // @[LoadUop.scala 80:62:@5613.4]
  wire [15:0] _T_76; // @[LoadUop.scala 80:88:@5614.4]
  wire [15:0] _T_77; // @[LoadUop.scala 80:88:@5615.4]
  wire [14:0] xsize; // @[LoadUop.scala 80:88:@5616.4]
  wire [31:0] _GEN_31; // @[LoadUop.scala 84:36:@5617.4]
  wire [1:0] _T_79; // @[LoadUop.scala 84:36:@5617.4]
  wire  dram_even; // @[LoadUop.scala 84:43:@5618.4]
  wire  sram_even; // @[LoadUop.scala 85:43:@5620.4]
  wire [15:0] _GEN_36; // @[LoadUop.scala 86:31:@5621.4]
  wire [1:0] _T_85; // @[LoadUop.scala 86:31:@5621.4]
  wire  sizeIsEven; // @[LoadUop.scala 86:38:@5622.4]
  reg [1:0] state; // @[LoadUop.scala 89:22:@5623.4]
  reg [31:0] _RAND_6;
  wire  _T_88; // @[Conditional.scala 37:30:@5624.4]
  wire  _T_89; // @[LoadUop.scala 96:20:@5628.8]
  wire [9:0] _T_92; // @[LoadUop.scala 100:24:@5634.10]
  wire [9:0] _T_93; // @[LoadUop.scala 100:24:@5635.10]
  wire [8:0] _T_94; // @[LoadUop.scala 100:24:@5636.10]
  wire [15:0] _T_95; // @[LoadUop.scala 101:25:@5638.10]
  wire [15:0] _T_96; // @[LoadUop.scala 101:25:@5639.10]
  wire [14:0] _T_97; // @[LoadUop.scala 101:25:@5640.10]
  wire [14:0] _GEN_0; // @[LoadUop.scala 96:28:@5629.8]
  wire [14:0] _GEN_1; // @[LoadUop.scala 96:28:@5629.8]
  wire [1:0] _GEN_2; // @[LoadUop.scala 94:22:@5626.6]
  wire [14:0] _GEN_3; // @[LoadUop.scala 94:22:@5626.6]
  wire [15:0] _GEN_4; // @[LoadUop.scala 94:22:@5626.6]
  wire  _T_98; // @[Conditional.scala 37:30:@5646.6]
  wire [1:0] _GEN_5; // @[LoadUop.scala 106:33:@5648.8]
  wire  _T_99; // @[Conditional.scala 37:30:@5653.8]
  wire  _T_100; // @[LoadUop.scala 112:19:@5656.12]
  wire  _T_102; // @[LoadUop.scala 113:21:@5658.14]
  wire [32:0] _T_103; // @[LoadUop.scala 116:28:@5663.16]
  wire [31:0] _T_104; // @[LoadUop.scala 116:28:@5664.16]
  wire  _T_105; // @[LoadUop.scala 117:23:@5666.16]
  wire [16:0] _T_111; // @[LoadUop.scala 125:28:@5678.18]
  wire [16:0] _T_112; // @[LoadUop.scala 125:28:@5679.18]
  wire [15:0] _T_113; // @[LoadUop.scala 125:28:@5680.18]
  wire [15:0] _GEN_7; // @[LoadUop.scala 117:31:@5667.16]
  wire [15:0] _GEN_8; // @[LoadUop.scala 117:31:@5667.16]
  wire [1:0] _GEN_9; // @[LoadUop.scala 113:30:@5659.14]
  wire [31:0] _GEN_10; // @[LoadUop.scala 113:30:@5659.14]
  wire [15:0] _GEN_11; // @[LoadUop.scala 113:30:@5659.14]
  wire [15:0] _GEN_12; // @[LoadUop.scala 113:30:@5659.14]
  wire [1:0] _GEN_13; // @[LoadUop.scala 112:29:@5657.12]
  wire [31:0] _GEN_14; // @[LoadUop.scala 112:29:@5657.12]
  wire [15:0] _GEN_15; // @[LoadUop.scala 112:29:@5657.12]
  wire [15:0] _GEN_16; // @[LoadUop.scala 112:29:@5657.12]
  wire [1:0] _GEN_17; // @[LoadUop.scala 111:34:@5655.10]
  wire [31:0] _GEN_18; // @[LoadUop.scala 111:34:@5655.10]
  wire [15:0] _GEN_19; // @[LoadUop.scala 111:34:@5655.10]
  wire [15:0] _GEN_20; // @[LoadUop.scala 111:34:@5655.10]
  wire [1:0] _GEN_21; // @[Conditional.scala 39:67:@5654.8]
  wire [31:0] _GEN_22; // @[Conditional.scala 39:67:@5654.8]
  wire [15:0] _GEN_23; // @[Conditional.scala 39:67:@5654.8]
  wire [15:0] _GEN_24; // @[Conditional.scala 39:67:@5654.8]
  wire [1:0] _GEN_25; // @[Conditional.scala 39:67:@5647.6]
  wire [31:0] _GEN_26; // @[Conditional.scala 39:67:@5647.6]
  wire [15:0] _GEN_27; // @[Conditional.scala 39:67:@5647.6]
  wire [15:0] _GEN_28; // @[Conditional.scala 39:67:@5647.6]
  wire [1:0] _GEN_29; // @[Conditional.scala 40:58:@5625.4]
  wire [15:0] _GEN_30; // @[Conditional.scala 40:58:@5625.4]
  wire [31:0] _GEN_32; // @[Conditional.scala 40:58:@5625.4]
  wire  _T_214; // @[LoadUop.scala 135:14:@5751.4]
  wire [33:0] _GEN_91; // @[LoadUop.scala 137:58:@5754.8]
  wire [33:0] _T_215; // @[LoadUop.scala 137:58:@5754.8]
  wire [33:0] _T_216; // @[LoadUop.scala 137:39:@5755.8]
  wire [33:0] _GEN_92; // @[LoadUop.scala 137:25:@5756.8]
  wire [33:0] _T_217; // @[LoadUop.scala 137:25:@5756.8]
  wire [34:0] _T_222; // @[LoadUop.scala 139:84:@5763.8]
  wire [34:0] _T_223; // @[LoadUop.scala 139:84:@5764.8]
  wire [33:0] _T_224; // @[LoadUop.scala 139:84:@5765.8]
  wire [33:0] _GEN_33; // @[LoadUop.scala 136:21:@5753.6]
  wire [33:0] _GEN_34; // @[LoadUop.scala 135:25:@5752.4]
  wire  _T_226; // @[LoadUop.scala 147:33:@5773.4]
  wire  _T_227; // @[LoadUop.scala 149:14:@5775.4]
  wire  _T_229; // @[Decoupled.scala 37:37:@5780.6]
  wire [8:0] _T_231; // @[LoadUop.scala 152:18:@5782.8]
  wire [7:0] _T_232; // @[LoadUop.scala 152:18:@5783.8]
  wire [7:0] _GEN_35; // @[LoadUop.scala 151:37:@5781.6]
  reg [9:0] waddr; // @[LoadUop.scala 155:18:@5786.4]
  reg [31:0] _RAND_7;
  wire [14:0] _T_235; // @[LoadUop.scala 157:30:@5789.6]
  wire [10:0] _T_238; // @[LoadUop.scala 159:20:@5795.8]
  wire [9:0] _T_239; // @[LoadUop.scala 159:20:@5796.8]
  wire [9:0] _GEN_37; // @[LoadUop.scala 158:37:@5794.6]
  wire [14:0] _GEN_38; // @[LoadUop.scala 156:25:@5788.4]
  reg  wmask_0; // @[LoadUop.scala 164:18:@5801.4]
  reg [31:0] _RAND_8;
  reg  wmask_1; // @[LoadUop.scala 164:18:@5801.4]
  reg [31:0] _RAND_9;
  wire  _T_297; // @[Decoupled.scala 37:37:@5815.8]
  wire  _T_299; // @[LoadUop.scala 170:22:@5817.10]
  wire  _GEN_40; // @[LoadUop.scala 170:31:@5818.10]
  wire [8:0] _T_350; // @[LoadUop.scala 176:27:@5844.12]
  wire [8:0] _T_351; // @[LoadUop.scala 176:27:@5845.12]
  wire [7:0] _T_352; // @[LoadUop.scala 176:27:@5846.12]
  wire  _T_353; // @[LoadUop.scala 176:18:@5847.12]
  wire  _T_356; // @[LoadUop.scala 176:34:@5849.12]
  wire  _GEN_42; // @[LoadUop.scala 176:53:@5850.12]
  wire  _GEN_43; // @[LoadUop.scala 175:39:@5843.10]
  wire  _GEN_44; // @[LoadUop.scala 175:39:@5843.10]
  wire  _GEN_45; // @[LoadUop.scala 169:38:@5816.8]
  wire  _GEN_46; // @[LoadUop.scala 169:38:@5816.8]
  wire  _GEN_47; // @[LoadUop.scala 167:22:@5803.6]
  wire  _GEN_48; // @[LoadUop.scala 167:22:@5803.6]
  wire  _T_436; // @[LoadUop.scala 186:23:@5894.10]
  wire  _T_439; // @[LoadUop.scala 186:48:@5896.10]
  wire  _GEN_50; // @[LoadUop.scala 186:67:@5897.10]
  wire  _GEN_52; // @[LoadUop.scala 185:39:@5889.8]
  wire  _GEN_53; // @[LoadUop.scala 183:32:@5876.6]
  wire  _GEN_54; // @[LoadUop.scala 183:32:@5876.6]
  wire [31:0] _T_509; // @[LoadUop.scala 194:40:@5924.4]
  wire [31:0] _T_510; // @[LoadUop.scala 194:40:@5926.4]
  wire  _T_512; // @[LoadUop.scala 195:18:@5930.4]
  wire  _T_513; // @[LoadUop.scala 195:30:@5931.4]
  wire  _T_538; // @[LoadUop.scala 197:24:@5943.6]
  wire  _T_539; // @[LoadUop.scala 197:36:@5944.6]
  wire [31:0] _GEN_57; // @[LoadUop.scala 197:50:@5945.6]
  reg  _T_579; // @[LoadUop.scala 206:31:@5965.4]
  reg [31:0] _RAND_10;
  wire [10:0] _GEN_39; // @[LoadUop.scala 208:30:@5968.4]
  wire [1:0] sIdx; // @[LoadUop.scala 208:30:@5968.4]
  wire [9:0] rIdx; // @[LoadUop.scala 209:30:@5969.4]
  wire  _GEN_72; // @[LoadUop.scala 210:25:@5972.4]
  wire [63:0] _T_599; // @[LoadUop.scala 211:23:@5978.4]
  wire [31:0] sWord_0; // @[LoadUop.scala 211:38:@5982.4]
  wire [31:0] sWord_1; // @[LoadUop.scala 211:38:@5984.4]
  wire  _T_625; // @[:@5986.4]
  wire [31:0] _GEN_76; // @[:@5989.4]
  wire  _T_633; // @[LoadUop.scala 217:34:@6000.4]
  wire  _T_635; // @[LoadUop.scala 217:57:@6002.4]
  reg [9:0] mem_0_memRead_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [9:0] mem_1_memRead_addr_pipe_0;
  reg [31:0] _RAND_12;
  assign mem_0_memRead_addr = mem_0_memRead_addr_pipe_0;
  assign mem_0_memRead_data = mem_0[mem_0_memRead_addr]; // @[LoadUop.scala 163:24:@5800.4]
  assign mem_0__T_564_data = _T_513 ? _T_510 : _T_509;
  assign mem_0__T_564_addr = waddr;
  assign mem_0__T_564_mask = wmask_0;
  assign mem_0__T_564_en = io_vme_rd_data_ready & io_vme_rd_data_valid;
  assign mem_1_memRead_addr = mem_1_memRead_addr_pipe_0;
  assign mem_1_memRead_data = mem_1[mem_1_memRead_addr]; // @[LoadUop.scala 163:24:@5800.4]
  assign mem_1__T_564_data = _T_513 ? _T_510 : _GEN_57;
  assign mem_1__T_564_addr = waddr;
  assign mem_1__T_564_mask = wmask_1;
  assign mem_1__T_564_en = io_vme_rd_data_ready & io_vme_rd_data_valid;
  assign dec_sram_offset = io_inst[24:9]; // @[LoadUop.scala 75:29:@5583.4]
  assign dec_dram_offset = io_inst[56:25]; // @[LoadUop.scala 75:29:@5585.4]
  assign dec_xsize = io_inst[95:80]; // @[LoadUop.scala 75:29:@5591.4]
  assign _T_67 = dec_xsize[15:1]; // @[LoadUop.scala 80:26:@5607.4]
  assign _T_68 = dec_xsize[0]; // @[LoadUop.scala 80:58:@5608.4]
  assign _GEN_89 = {{14'd0}, _T_68}; // @[LoadUop.scala 80:47:@5609.4]
  assign _T_69 = _T_67 + _GEN_89; // @[LoadUop.scala 80:47:@5609.4]
  assign _T_70 = _T_67 + _GEN_89; // @[LoadUop.scala 80:47:@5610.4]
  assign _GEN_6 = dec_sram_offset % 16'h2; // @[LoadUop.scala 80:81:@5611.4]
  assign _T_72 = _GEN_6[1:0]; // @[LoadUop.scala 80:81:@5611.4]
  assign _GEN_90 = {{13'd0}, _T_72}; // @[LoadUop.scala 80:62:@5612.4]
  assign _T_73 = _T_70 + _GEN_90; // @[LoadUop.scala 80:62:@5612.4]
  assign _T_74 = _T_70 + _GEN_90; // @[LoadUop.scala 80:62:@5613.4]
  assign _T_76 = _T_74 - 15'h1; // @[LoadUop.scala 80:88:@5614.4]
  assign _T_77 = $unsigned(_T_76); // @[LoadUop.scala 80:88:@5615.4]
  assign xsize = _T_77[14:0]; // @[LoadUop.scala 80:88:@5616.4]
  assign _GEN_31 = dec_dram_offset % 32'h2; // @[LoadUop.scala 84:36:@5617.4]
  assign _T_79 = _GEN_31[1:0]; // @[LoadUop.scala 84:36:@5617.4]
  assign dram_even = _T_79 == 2'h0; // @[LoadUop.scala 84:43:@5618.4]
  assign sram_even = _T_72 == 2'h0; // @[LoadUop.scala 85:43:@5620.4]
  assign _GEN_36 = dec_xsize % 16'h2; // @[LoadUop.scala 86:31:@5621.4]
  assign _T_85 = _GEN_36[1:0]; // @[LoadUop.scala 86:31:@5621.4]
  assign sizeIsEven = _T_85 == 2'h0; // @[LoadUop.scala 86:38:@5622.4]
  assign _T_88 = 2'h0 == state; // @[Conditional.scala 37:30:@5624.4]
  assign _T_89 = xsize < 15'h100; // @[LoadUop.scala 96:20:@5628.8]
  assign _T_92 = 9'h100 - 9'h1; // @[LoadUop.scala 100:24:@5634.10]
  assign _T_93 = $unsigned(_T_92); // @[LoadUop.scala 100:24:@5635.10]
  assign _T_94 = _T_93[8:0]; // @[LoadUop.scala 100:24:@5636.10]
  assign _T_95 = xsize - 15'h100; // @[LoadUop.scala 101:25:@5638.10]
  assign _T_96 = $unsigned(_T_95); // @[LoadUop.scala 101:25:@5639.10]
  assign _T_97 = _T_96[14:0]; // @[LoadUop.scala 101:25:@5640.10]
  assign _GEN_0 = _T_89 ? xsize : {{6'd0}, _T_94}; // @[LoadUop.scala 96:28:@5629.8]
  assign _GEN_1 = _T_89 ? 15'h0 : _T_97; // @[LoadUop.scala 96:28:@5629.8]
  assign _GEN_2 = io_start ? 2'h1 : state; // @[LoadUop.scala 94:22:@5626.6]
  assign _GEN_3 = io_start ? _GEN_0 : {{7'd0}, xlen}; // @[LoadUop.scala 94:22:@5626.6]
  assign _GEN_4 = io_start ? {{1'd0}, _GEN_1} : xrem; // @[LoadUop.scala 94:22:@5626.6]
  assign _T_98 = 2'h1 == state; // @[Conditional.scala 37:30:@5646.6]
  assign _GEN_5 = io_vme_rd_cmd_ready ? 2'h2 : state; // @[LoadUop.scala 106:33:@5648.8]
  assign _T_99 = 2'h2 == state; // @[Conditional.scala 37:30:@5653.8]
  assign _T_100 = xcnt == xlen; // @[LoadUop.scala 112:19:@5656.12]
  assign _T_102 = xrem == 16'h0; // @[LoadUop.scala 113:21:@5658.14]
  assign _T_103 = raddr + 32'h800; // @[LoadUop.scala 116:28:@5663.16]
  assign _T_104 = raddr + 32'h800; // @[LoadUop.scala 116:28:@5664.16]
  assign _T_105 = xrem < 16'h100; // @[LoadUop.scala 117:23:@5666.16]
  assign _T_111 = xrem - 16'h100; // @[LoadUop.scala 125:28:@5678.18]
  assign _T_112 = $unsigned(_T_111); // @[LoadUop.scala 125:28:@5679.18]
  assign _T_113 = _T_112[15:0]; // @[LoadUop.scala 125:28:@5680.18]
  assign _GEN_7 = _T_105 ? xrem : {{7'd0}, _T_94}; // @[LoadUop.scala 117:31:@5667.16]
  assign _GEN_8 = _T_105 ? 16'h0 : _T_113; // @[LoadUop.scala 117:31:@5667.16]
  assign _GEN_9 = _T_102 ? 2'h0 : 2'h1; // @[LoadUop.scala 113:30:@5659.14]
  assign _GEN_10 = _T_102 ? raddr : _T_104; // @[LoadUop.scala 113:30:@5659.14]
  assign _GEN_11 = _T_102 ? {{8'd0}, xlen} : _GEN_7; // @[LoadUop.scala 113:30:@5659.14]
  assign _GEN_12 = _T_102 ? xrem : _GEN_8; // @[LoadUop.scala 113:30:@5659.14]
  assign _GEN_13 = _T_100 ? _GEN_9 : state; // @[LoadUop.scala 112:29:@5657.12]
  assign _GEN_14 = _T_100 ? _GEN_10 : raddr; // @[LoadUop.scala 112:29:@5657.12]
  assign _GEN_15 = _T_100 ? _GEN_11 : {{8'd0}, xlen}; // @[LoadUop.scala 112:29:@5657.12]
  assign _GEN_16 = _T_100 ? _GEN_12 : xrem; // @[LoadUop.scala 112:29:@5657.12]
  assign _GEN_17 = io_vme_rd_data_valid ? _GEN_13 : state; // @[LoadUop.scala 111:34:@5655.10]
  assign _GEN_18 = io_vme_rd_data_valid ? _GEN_14 : raddr; // @[LoadUop.scala 111:34:@5655.10]
  assign _GEN_19 = io_vme_rd_data_valid ? _GEN_15 : {{8'd0}, xlen}; // @[LoadUop.scala 111:34:@5655.10]
  assign _GEN_20 = io_vme_rd_data_valid ? _GEN_16 : xrem; // @[LoadUop.scala 111:34:@5655.10]
  assign _GEN_21 = _T_99 ? _GEN_17 : state; // @[Conditional.scala 39:67:@5654.8]
  assign _GEN_22 = _T_99 ? _GEN_18 : raddr; // @[Conditional.scala 39:67:@5654.8]
  assign _GEN_23 = _T_99 ? _GEN_19 : {{8'd0}, xlen}; // @[Conditional.scala 39:67:@5654.8]
  assign _GEN_24 = _T_99 ? _GEN_20 : xrem; // @[Conditional.scala 39:67:@5654.8]
  assign _GEN_25 = _T_98 ? _GEN_5 : _GEN_21; // @[Conditional.scala 39:67:@5647.6]
  assign _GEN_26 = _T_98 ? raddr : _GEN_22; // @[Conditional.scala 39:67:@5647.6]
  assign _GEN_27 = _T_98 ? {{8'd0}, xlen} : _GEN_23; // @[Conditional.scala 39:67:@5647.6]
  assign _GEN_28 = _T_98 ? xrem : _GEN_24; // @[Conditional.scala 39:67:@5647.6]
  assign _GEN_29 = _T_88 ? _GEN_2 : _GEN_25; // @[Conditional.scala 40:58:@5625.4]
  assign _GEN_30 = _T_88 ? {{1'd0}, _GEN_3} : _GEN_27; // @[Conditional.scala 40:58:@5625.4]
  assign _GEN_32 = _T_88 ? raddr : _GEN_26; // @[Conditional.scala 40:58:@5625.4]
  assign _T_214 = state == 2'h0; // @[LoadUop.scala 135:14:@5751.4]
  assign _GEN_91 = {{2'd0}, dec_dram_offset}; // @[LoadUop.scala 137:58:@5754.8]
  assign _T_215 = _GEN_91 << 2; // @[LoadUop.scala 137:58:@5754.8]
  assign _T_216 = 34'hffffffff & _T_215; // @[LoadUop.scala 137:39:@5755.8]
  assign _GEN_92 = {{2'd0}, io_baddr}; // @[LoadUop.scala 137:25:@5756.8]
  assign _T_217 = _GEN_92 | _T_216; // @[LoadUop.scala 137:25:@5756.8]
  assign _T_222 = _T_217 - 34'h4; // @[LoadUop.scala 139:84:@5763.8]
  assign _T_223 = $unsigned(_T_222); // @[LoadUop.scala 139:84:@5764.8]
  assign _T_224 = _T_223[33:0]; // @[LoadUop.scala 139:84:@5765.8]
  assign _GEN_33 = dram_even ? _T_217 : _T_224; // @[LoadUop.scala 136:21:@5753.6]
  assign _GEN_34 = _T_214 ? _GEN_33 : {{2'd0}, _GEN_32}; // @[LoadUop.scala 135:25:@5752.4]
  assign _T_226 = state == 2'h2; // @[LoadUop.scala 147:33:@5773.4]
  assign _T_227 = state != 2'h2; // @[LoadUop.scala 149:14:@5775.4]
  assign _T_229 = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[Decoupled.scala 37:37:@5780.6]
  assign _T_231 = xcnt + 8'h1; // @[LoadUop.scala 152:18:@5782.8]
  assign _T_232 = xcnt + 8'h1; // @[LoadUop.scala 152:18:@5783.8]
  assign _GEN_35 = _T_229 ? _T_232 : xcnt; // @[LoadUop.scala 151:37:@5781.6]
  assign _T_235 = dec_sram_offset[15:1]; // @[LoadUop.scala 157:30:@5789.6]
  assign _T_238 = waddr + 10'h1; // @[LoadUop.scala 159:20:@5795.8]
  assign _T_239 = waddr + 10'h1; // @[LoadUop.scala 159:20:@5796.8]
  assign _GEN_37 = _T_229 ? _T_239 : waddr; // @[LoadUop.scala 158:37:@5794.6]
  assign _GEN_38 = _T_214 ? _T_235 : {{5'd0}, _GEN_37}; // @[LoadUop.scala 156:25:@5788.4]
  assign _T_297 = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[Decoupled.scala 37:37:@5815.8]
  assign _T_299 = dec_xsize == 16'h1; // @[LoadUop.scala 170:22:@5817.10]
  assign _GEN_40 = _T_299 ? 1'h0 : 1'h1; // @[LoadUop.scala 170:31:@5818.10]
  assign _T_350 = xlen - 8'h1; // @[LoadUop.scala 176:27:@5844.12]
  assign _T_351 = $unsigned(_T_350); // @[LoadUop.scala 176:27:@5845.12]
  assign _T_352 = _T_351[7:0]; // @[LoadUop.scala 176:27:@5846.12]
  assign _T_353 = xcnt == _T_352; // @[LoadUop.scala 176:18:@5847.12]
  assign _T_356 = _T_353 & _T_102; // @[LoadUop.scala 176:34:@5849.12]
  assign _GEN_42 = _T_356 ? 1'h0 : 1'h1; // @[LoadUop.scala 176:53:@5850.12]
  assign _GEN_43 = _T_229 ? 1'h1 : wmask_0; // @[LoadUop.scala 175:39:@5843.10]
  assign _GEN_44 = _T_229 ? _GEN_42 : wmask_1; // @[LoadUop.scala 175:39:@5843.10]
  assign _GEN_45 = _T_297 ? 1'h1 : _GEN_43; // @[LoadUop.scala 169:38:@5816.8]
  assign _GEN_46 = _T_297 ? _GEN_40 : _GEN_44; // @[LoadUop.scala 169:38:@5816.8]
  assign _GEN_47 = sizeIsEven ? 1'h1 : _GEN_45; // @[LoadUop.scala 167:22:@5803.6]
  assign _GEN_48 = sizeIsEven ? 1'h1 : _GEN_46; // @[LoadUop.scala 167:22:@5803.6]
  assign _T_436 = sizeIsEven & _T_353; // @[LoadUop.scala 186:23:@5894.10]
  assign _T_439 = _T_436 & _T_102; // @[LoadUop.scala 186:48:@5896.10]
  assign _GEN_50 = _T_439 ? 1'h0 : 1'h1; // @[LoadUop.scala 186:67:@5897.10]
  assign _GEN_52 = _T_229 ? _GEN_50 : wmask_1; // @[LoadUop.scala 185:39:@5889.8]
  assign _GEN_53 = _T_297 ? 1'h0 : _GEN_43; // @[LoadUop.scala 183:32:@5876.6]
  assign _GEN_54 = _T_297 ? 1'h1 : _GEN_52; // @[LoadUop.scala 183:32:@5876.6]
  assign _T_509 = io_vme_rd_data_bits[31:0]; // @[LoadUop.scala 194:40:@5924.4]
  assign _T_510 = io_vme_rd_data_bits[63:32]; // @[LoadUop.scala 194:40:@5926.4]
  assign _T_512 = dram_even == 1'h0; // @[LoadUop.scala 195:18:@5930.4]
  assign _T_513 = _T_512 & sram_even; // @[LoadUop.scala 195:30:@5931.4]
  assign _T_538 = sram_even == 1'h0; // @[LoadUop.scala 197:24:@5943.6]
  assign _T_539 = _T_538 & dram_even; // @[LoadUop.scala 197:36:@5944.6]
  assign _GEN_57 = _T_539 ? _T_509 : _T_510; // @[LoadUop.scala 197:50:@5945.6]
  assign _GEN_39 = io_uop_idx_bits % 11'h2; // @[LoadUop.scala 208:30:@5968.4]
  assign sIdx = _GEN_39[1:0]; // @[LoadUop.scala 208:30:@5968.4]
  assign rIdx = io_uop_idx_bits[10:1]; // @[LoadUop.scala 209:30:@5969.4]
  assign _GEN_72 = io_uop_idx_valid; // @[LoadUop.scala 210:25:@5972.4]
  assign _T_599 = {mem_1_memRead_data,mem_0_memRead_data}; // @[LoadUop.scala 211:23:@5978.4]
  assign sWord_0 = _T_599[31:0]; // @[LoadUop.scala 211:38:@5982.4]
  assign sWord_1 = _T_599[63:32]; // @[LoadUop.scala 211:38:@5984.4]
  assign _T_625 = sIdx[0]; // @[:@5986.4]
  assign _GEN_76 = _T_625 ? sWord_1 : sWord_0; // @[:@5989.4]
  assign _T_633 = _T_226 & io_vme_rd_data_valid; // @[LoadUop.scala 217:34:@6000.4]
  assign _T_635 = _T_633 & _T_100; // @[LoadUop.scala 217:57:@6002.4]
  assign io_done = _T_635 & _T_102; // @[LoadUop.scala 217:11:@6005.4]
  assign io_vme_rd_cmd_valid = state == 2'h1; // @[LoadUop.scala 143:23:@5770.4]
  assign io_vme_rd_cmd_bits_addr = raddr; // @[LoadUop.scala 144:27:@5771.4]
  assign io_vme_rd_cmd_bits_len = xlen; // @[LoadUop.scala 145:26:@5772.4]
  assign io_vme_rd_data_ready = state == 2'h2; // @[LoadUop.scala 147:24:@5774.4]
  assign io_uop_data_valid = _T_579; // @[LoadUop.scala 206:21:@5967.4]
  assign io_uop_data_bits_u2 = _GEN_76[31:22]; // @[LoadUop.scala 214:20:@5998.4]
  assign io_uop_data_bits_u1 = _GEN_76[21:11]; // @[LoadUop.scala 214:20:@5997.4]
  assign io_uop_data_bits_u0 = _GEN_76[10:0]; // @[LoadUop.scala 214:20:@5996.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem_0[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem_1[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  raddr = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  xcnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xlen = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  xrem = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  waddr = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wmask_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wmask_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_579 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_0_memRead_addr_pipe_0 = _RAND_11[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mem_1_memRead_addr_pipe_0 = _RAND_12[9:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem_0__T_564_en & mem_0__T_564_mask) begin
      mem_0[mem_0__T_564_addr] <= mem_0__T_564_data; // @[LoadUop.scala 163:24:@5800.4]
    end
    if(mem_1__T_564_en & mem_1__T_564_mask) begin
      mem_1[mem_1__T_564_addr] <= mem_1__T_564_data; // @[LoadUop.scala 163:24:@5800.4]
    end
    raddr <= _GEN_34[31:0];
    if (_T_227) begin
      xcnt <= 8'h0;
    end else begin
      if (_T_229) begin
        xcnt <= _T_232;
      end
    end
    xlen <= _GEN_30[7:0];
    if (_T_88) begin
      if (io_start) begin
        xrem <= {{1'd0}, _GEN_1};
      end
    end else begin
      if (!(_T_98)) begin
        if (_T_99) begin
          if (io_vme_rd_data_valid) begin
            if (_T_100) begin
              if (!(_T_102)) begin
                if (_T_105) begin
                  xrem <= 16'h0;
                end else begin
                  xrem <= _T_113;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_88) begin
        if (io_start) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_98) begin
          if (io_vme_rd_cmd_ready) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_99) begin
            if (io_vme_rd_data_valid) begin
              if (_T_100) begin
                if (_T_102) begin
                  state <= 2'h0;
                end else begin
                  state <= 2'h1;
                end
              end
            end
          end
        end
      end
    end
    waddr <= _GEN_38[9:0];
    if (sram_even) begin
      if (sizeIsEven) begin
        wmask_0 <= 1'h1;
      end else begin
        if (_T_297) begin
          wmask_0 <= 1'h1;
        end else begin
          if (_T_229) begin
            wmask_0 <= 1'h1;
          end
        end
      end
    end else begin
      if (_T_297) begin
        wmask_0 <= 1'h0;
      end else begin
        if (_T_229) begin
          wmask_0 <= 1'h1;
        end
      end
    end
    if (sram_even) begin
      if (sizeIsEven) begin
        wmask_1 <= 1'h1;
      end else begin
        if (_T_297) begin
          if (_T_299) begin
            wmask_1 <= 1'h0;
          end else begin
            wmask_1 <= 1'h1;
          end
        end else begin
          if (_T_229) begin
            if (_T_356) begin
              wmask_1 <= 1'h0;
            end else begin
              wmask_1 <= 1'h1;
            end
          end
        end
      end
    end else begin
      if (_T_297) begin
        wmask_1 <= 1'h1;
      end else begin
        if (_T_229) begin
          if (_T_439) begin
            wmask_1 <= 1'h0;
          end else begin
            wmask_1 <= 1'h1;
          end
        end
      end
    end
    _T_579 <= io_uop_idx_valid;
    if (_GEN_72) begin
      mem_0_memRead_addr_pipe_0 <= rIdx;
    end
    if (_GEN_72) begin
      mem_1_memRead_addr_pipe_0 <= rIdx;
    end
  end
endmodule
module TensorDataCtrl_2( // @[:@6007.2]
  input          clock, // @[:@6008.4]
  input          io_start, // @[:@6010.4]
  output         io_done, // @[:@6010.4]
  input  [127:0] io_inst, // @[:@6010.4]
  input  [31:0]  io_baddr, // @[:@6010.4]
  input          io_xinit, // @[:@6010.4]
  input          io_xupdate, // @[:@6010.4]
  input          io_yupdate, // @[:@6010.4]
  output         io_stride, // @[:@6010.4]
  output         io_split, // @[:@6010.4]
  output [31:0]  io_addr, // @[:@6010.4]
  output [7:0]   io_len // @[:@6010.4]
);
  wire [31:0] dec_dram_offset; // @[TensorUtil.scala 251:29:@6029.4]
  wire [15:0] dec_ysize; // @[TensorUtil.scala 251:29:@6033.4]
  wire [15:0] dec_xsize; // @[TensorUtil.scala 251:29:@6035.4]
  wire [15:0] dec_xstride; // @[TensorUtil.scala 251:29:@6037.4]
  reg [31:0] caddr; // @[TensorUtil.scala 253:18:@6047.4]
  reg [31:0] _RAND_0;
  reg [31:0] baddr; // @[TensorUtil.scala 254:18:@6048.4]
  reg [31:0] _RAND_1;
  reg [7:0] len; // @[TensorUtil.scala 255:16:@6049.4]
  reg [31:0] _RAND_2;
  reg [7:0] xcnt; // @[TensorUtil.scala 267:17:@6114.4]
  reg [31:0] _RAND_3;
  reg [15:0] xrem; // @[TensorUtil.scala 268:17:@6115.4]
  reg [31:0] _RAND_4;
  wire [18:0] _GEN_27; // @[TensorUtil.scala 269:26:@6116.4]
  wire [18:0] _T_154; // @[TensorUtil.scala 269:26:@6116.4]
  wire [19:0] _T_156; // @[TensorUtil.scala 269:51:@6117.4]
  wire [19:0] _T_157; // @[TensorUtil.scala 269:51:@6118.4]
  wire [18:0] xsize; // @[TensorUtil.scala 269:51:@6119.4]
  reg [15:0] ycnt; // @[TensorUtil.scala 271:17:@6120.4]
  reg [31:0] _RAND_5;
  reg [31:0] xfer_bytes; // @[TensorUtil.scala 273:23:@6121.4]
  reg [31:0] _RAND_6;
  wire [21:0] _GEN_28; // @[TensorUtil.scala 275:35:@6122.4]
  wire [21:0] xstride_bytes; // @[TensorUtil.scala 275:35:@6122.4]
  wire [37:0] _GEN_29; // @[TensorUtil.scala 277:66:@6123.4]
  wire [37:0] _T_160; // @[TensorUtil.scala 277:66:@6123.4]
  wire [37:0] _T_161; // @[TensorUtil.scala 277:47:@6124.4]
  wire [37:0] _GEN_30; // @[TensorUtil.scala 277:33:@6125.4]
  wire [37:0] xfer_init_addr; // @[TensorUtil.scala 277:33:@6125.4]
  wire [32:0] _T_162; // @[TensorUtil.scala 278:31:@6126.4]
  wire [31:0] xfer_split_addr; // @[TensorUtil.scala 278:31:@6127.4]
  wire [31:0] _GEN_31; // @[TensorUtil.scala 279:32:@6128.4]
  wire [32:0] _T_163; // @[TensorUtil.scala 279:32:@6128.4]
  wire [31:0] xfer_stride_addr; // @[TensorUtil.scala 279:32:@6129.4]
  wire [37:0] _GEN_12; // @[TensorUtil.scala 281:55:@6130.4]
  wire [11:0] _T_164; // @[TensorUtil.scala 281:55:@6130.4]
  wire [12:0] _T_165; // @[TensorUtil.scala 281:38:@6131.4]
  wire [12:0] _T_166; // @[TensorUtil.scala 281:38:@6132.4]
  wire [11:0] xfer_init_bytes; // @[TensorUtil.scala 281:38:@6133.4]
  wire [8:0] xfer_init_pulses; // @[TensorUtil.scala 282:43:@6134.4]
  wire [31:0] _GEN_16; // @[TensorUtil.scala 283:56:@6135.4]
  wire [11:0] _T_167; // @[TensorUtil.scala 283:56:@6135.4]
  wire [12:0] _T_168; // @[TensorUtil.scala 283:38:@6136.4]
  wire [12:0] _T_169; // @[TensorUtil.scala 283:38:@6137.4]
  wire [11:0] xfer_split_bytes; // @[TensorUtil.scala 283:38:@6138.4]
  wire [8:0] xfer_split_pulses; // @[TensorUtil.scala 284:44:@6139.4]
  wire [31:0] _GEN_18; // @[TensorUtil.scala 285:57:@6140.4]
  wire [11:0] _T_170; // @[TensorUtil.scala 285:57:@6140.4]
  wire [12:0] _T_171; // @[TensorUtil.scala 285:38:@6141.4]
  wire [12:0] _T_172; // @[TensorUtil.scala 285:38:@6142.4]
  wire [11:0] xfer_stride_bytes; // @[TensorUtil.scala 285:38:@6143.4]
  wire [8:0] xfer_stride_pulses; // @[TensorUtil.scala 286:45:@6144.4]
  wire  _T_173; // @[TensorUtil.scala 288:21:@6145.4]
  wire  _T_175; // @[TensorUtil.scala 289:10:@6146.4]
  wire  _T_176; // @[TensorUtil.scala 288:29:@6147.4]
  wire [16:0] _T_178; // @[TensorUtil.scala 290:24:@6148.4]
  wire [16:0] _T_179; // @[TensorUtil.scala 290:24:@6149.4]
  wire [15:0] _T_180; // @[TensorUtil.scala 290:24:@6150.4]
  wire  _T_181; // @[TensorUtil.scala 290:10:@6151.4]
  wire  stride; // @[TensorUtil.scala 289:18:@6152.4]
  wire  _T_184; // @[TensorUtil.scala 292:35:@6154.4]
  wire  split; // @[TensorUtil.scala 292:28:@6155.4]
  wire [18:0] _GEN_32; // @[TensorUtil.scala 296:16:@6158.6]
  wire  _T_185; // @[TensorUtil.scala 296:16:@6158.6]
  wire [9:0] _T_188; // @[TensorUtil.scala 300:31:@6164.8]
  wire [9:0] _T_189; // @[TensorUtil.scala 300:31:@6165.8]
  wire [8:0] _T_190; // @[TensorUtil.scala 300:31:@6166.8]
  wire [19:0] _T_191; // @[TensorUtil.scala 301:21:@6168.8]
  wire [19:0] _T_192; // @[TensorUtil.scala 301:21:@6169.8]
  wire [18:0] _T_193; // @[TensorUtil.scala 301:21:@6170.8]
  wire [18:0] _GEN_0; // @[TensorUtil.scala 296:36:@6159.6]
  wire [18:0] _GEN_1; // @[TensorUtil.scala 296:36:@6159.6]
  wire  _T_194; // @[TensorUtil.scala 303:25:@6175.6]
  wire [18:0] _GEN_34; // @[TensorUtil.scala 305:16:@6178.8]
  wire  _T_195; // @[TensorUtil.scala 305:16:@6178.8]
  wire [9:0] _T_198; // @[TensorUtil.scala 309:33:@6184.10]
  wire [9:0] _T_199; // @[TensorUtil.scala 309:33:@6185.10]
  wire [8:0] _T_200; // @[TensorUtil.scala 309:33:@6186.10]
  wire [19:0] _T_201; // @[TensorUtil.scala 310:21:@6188.10]
  wire [19:0] _T_202; // @[TensorUtil.scala 310:21:@6189.10]
  wire [18:0] _T_203; // @[TensorUtil.scala 310:21:@6190.10]
  wire [18:0] _GEN_2; // @[TensorUtil.scala 305:38:@6179.8]
  wire [18:0] _GEN_3; // @[TensorUtil.scala 305:38:@6179.8]
  wire  _T_204; // @[TensorUtil.scala 312:25:@6195.8]
  wire [15:0] _GEN_36; // @[TensorUtil.scala 314:15:@6198.10]
  wire  _T_205; // @[TensorUtil.scala 314:15:@6198.10]
  wire [9:0] _T_208; // @[TensorUtil.scala 318:32:@6204.12]
  wire [9:0] _T_209; // @[TensorUtil.scala 318:32:@6205.12]
  wire [8:0] _T_210; // @[TensorUtil.scala 318:32:@6206.12]
  wire [16:0] _T_211; // @[TensorUtil.scala 319:20:@6208.12]
  wire [16:0] _T_212; // @[TensorUtil.scala 319:20:@6209.12]
  wire [15:0] _T_213; // @[TensorUtil.scala 319:20:@6210.12]
  wire [15:0] _GEN_4; // @[TensorUtil.scala 314:36:@6199.10]
  wire [15:0] _GEN_5; // @[TensorUtil.scala 314:36:@6199.10]
  wire [31:0] _GEN_6; // @[TensorUtil.scala 312:35:@6196.8]
  wire [15:0] _GEN_7; // @[TensorUtil.scala 312:35:@6196.8]
  wire [15:0] _GEN_8; // @[TensorUtil.scala 312:35:@6196.8]
  wire [31:0] _GEN_9; // @[TensorUtil.scala 303:36:@6176.6]
  wire [18:0] _GEN_10; // @[TensorUtil.scala 303:36:@6176.6]
  wire [18:0] _GEN_11; // @[TensorUtil.scala 303:36:@6176.6]
  wire [18:0] _GEN_13; // @[TensorUtil.scala 294:18:@6156.4]
  wire [18:0] _GEN_14; // @[TensorUtil.scala 294:18:@6156.4]
  wire [8:0] _T_216; // @[TensorUtil.scala 326:18:@6219.8]
  wire [7:0] _T_217; // @[TensorUtil.scala 326:18:@6220.8]
  wire [7:0] _GEN_15; // @[TensorUtil.scala 325:26:@6218.6]
  wire  _T_219; // @[TensorUtil.scala 331:25:@6227.6]
  wire [16:0] _T_221; // @[TensorUtil.scala 332:18:@6229.8]
  wire [15:0] _T_222; // @[TensorUtil.scala 332:18:@6230.8]
  wire [15:0] _GEN_17; // @[TensorUtil.scala 331:36:@6228.6]
  wire [31:0] _GEN_19; // @[TensorUtil.scala 341:24:@6243.10]
  wire [31:0] _GEN_20; // @[TensorUtil.scala 341:24:@6243.10]
  wire [31:0] _GEN_21; // @[TensorUtil.scala 339:17:@6239.8]
  wire [31:0] _GEN_22; // @[TensorUtil.scala 339:17:@6239.8]
  wire [31:0] _GEN_23; // @[TensorUtil.scala 338:26:@6238.6]
  wire [31:0] _GEN_24; // @[TensorUtil.scala 338:26:@6238.6]
  wire [37:0] _GEN_25; // @[TensorUtil.scala 335:18:@6233.4]
  wire [37:0] _GEN_26; // @[TensorUtil.scala 335:18:@6233.4]
  wire  _T_232; // @[TensorUtil.scala 354:10:@6260.4]
  assign dec_dram_offset = io_inst[56:25]; // @[TensorUtil.scala 251:29:@6029.4]
  assign dec_ysize = io_inst[79:64]; // @[TensorUtil.scala 251:29:@6033.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 251:29:@6035.4]
  assign dec_xstride = io_inst[111:96]; // @[TensorUtil.scala 251:29:@6037.4]
  assign _GEN_27 = {{3'd0}, dec_xsize}; // @[TensorUtil.scala 269:26:@6116.4]
  assign _T_154 = _GEN_27 << 3; // @[TensorUtil.scala 269:26:@6116.4]
  assign _T_156 = _T_154 - 19'h1; // @[TensorUtil.scala 269:51:@6117.4]
  assign _T_157 = $unsigned(_T_156); // @[TensorUtil.scala 269:51:@6118.4]
  assign xsize = _T_157[18:0]; // @[TensorUtil.scala 269:51:@6119.4]
  assign _GEN_28 = {{6'd0}, dec_xstride}; // @[TensorUtil.scala 275:35:@6122.4]
  assign xstride_bytes = _GEN_28 << 6; // @[TensorUtil.scala 275:35:@6122.4]
  assign _GEN_29 = {{6'd0}, dec_dram_offset}; // @[TensorUtil.scala 277:66:@6123.4]
  assign _T_160 = _GEN_29 << 6; // @[TensorUtil.scala 277:66:@6123.4]
  assign _T_161 = 38'hffffffff & _T_160; // @[TensorUtil.scala 277:47:@6124.4]
  assign _GEN_30 = {{6'd0}, io_baddr}; // @[TensorUtil.scala 277:33:@6125.4]
  assign xfer_init_addr = _GEN_30 | _T_161; // @[TensorUtil.scala 277:33:@6125.4]
  assign _T_162 = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@6126.4]
  assign xfer_split_addr = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@6127.4]
  assign _GEN_31 = {{10'd0}, xstride_bytes}; // @[TensorUtil.scala 279:32:@6128.4]
  assign _T_163 = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@6128.4]
  assign xfer_stride_addr = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@6129.4]
  assign _GEN_12 = xfer_init_addr % 38'h800; // @[TensorUtil.scala 281:55:@6130.4]
  assign _T_164 = _GEN_12[11:0]; // @[TensorUtil.scala 281:55:@6130.4]
  assign _T_165 = 12'h800 - _T_164; // @[TensorUtil.scala 281:38:@6131.4]
  assign _T_166 = $unsigned(_T_165); // @[TensorUtil.scala 281:38:@6132.4]
  assign xfer_init_bytes = _T_166[11:0]; // @[TensorUtil.scala 281:38:@6133.4]
  assign xfer_init_pulses = xfer_init_bytes[11:3]; // @[TensorUtil.scala 282:43:@6134.4]
  assign _GEN_16 = xfer_split_addr % 32'h800; // @[TensorUtil.scala 283:56:@6135.4]
  assign _T_167 = _GEN_16[11:0]; // @[TensorUtil.scala 283:56:@6135.4]
  assign _T_168 = 12'h800 - _T_167; // @[TensorUtil.scala 283:38:@6136.4]
  assign _T_169 = $unsigned(_T_168); // @[TensorUtil.scala 283:38:@6137.4]
  assign xfer_split_bytes = _T_169[11:0]; // @[TensorUtil.scala 283:38:@6138.4]
  assign xfer_split_pulses = xfer_split_bytes[11:3]; // @[TensorUtil.scala 284:44:@6139.4]
  assign _GEN_18 = xfer_stride_addr % 32'h800; // @[TensorUtil.scala 285:57:@6140.4]
  assign _T_170 = _GEN_18[11:0]; // @[TensorUtil.scala 285:57:@6140.4]
  assign _T_171 = 12'h800 - _T_170; // @[TensorUtil.scala 285:38:@6141.4]
  assign _T_172 = $unsigned(_T_171); // @[TensorUtil.scala 285:38:@6142.4]
  assign xfer_stride_bytes = _T_172[11:0]; // @[TensorUtil.scala 285:38:@6143.4]
  assign xfer_stride_pulses = xfer_stride_bytes[11:3]; // @[TensorUtil.scala 286:45:@6144.4]
  assign _T_173 = xcnt == len; // @[TensorUtil.scala 288:21:@6145.4]
  assign _T_175 = xrem == 16'h0; // @[TensorUtil.scala 289:10:@6146.4]
  assign _T_176 = _T_173 & _T_175; // @[TensorUtil.scala 288:29:@6147.4]
  assign _T_178 = dec_ysize - 16'h1; // @[TensorUtil.scala 290:24:@6148.4]
  assign _T_179 = $unsigned(_T_178); // @[TensorUtil.scala 290:24:@6149.4]
  assign _T_180 = _T_179[15:0]; // @[TensorUtil.scala 290:24:@6150.4]
  assign _T_181 = ycnt != _T_180; // @[TensorUtil.scala 290:10:@6151.4]
  assign stride = _T_176 & _T_181; // @[TensorUtil.scala 289:18:@6152.4]
  assign _T_184 = xrem != 16'h0; // @[TensorUtil.scala 292:35:@6154.4]
  assign split = _T_173 & _T_184; // @[TensorUtil.scala 292:28:@6155.4]
  assign _GEN_32 = {{10'd0}, xfer_init_pulses}; // @[TensorUtil.scala 296:16:@6158.6]
  assign _T_185 = xsize < _GEN_32; // @[TensorUtil.scala 296:16:@6158.6]
  assign _T_188 = xfer_init_pulses - 9'h1; // @[TensorUtil.scala 300:31:@6164.8]
  assign _T_189 = $unsigned(_T_188); // @[TensorUtil.scala 300:31:@6165.8]
  assign _T_190 = _T_189[8:0]; // @[TensorUtil.scala 300:31:@6166.8]
  assign _T_191 = xsize - _GEN_32; // @[TensorUtil.scala 301:21:@6168.8]
  assign _T_192 = $unsigned(_T_191); // @[TensorUtil.scala 301:21:@6169.8]
  assign _T_193 = _T_192[18:0]; // @[TensorUtil.scala 301:21:@6170.8]
  assign _GEN_0 = _T_185 ? xsize : {{10'd0}, _T_190}; // @[TensorUtil.scala 296:36:@6159.6]
  assign _GEN_1 = _T_185 ? 19'h0 : _T_193; // @[TensorUtil.scala 296:36:@6159.6]
  assign _T_194 = io_xupdate & stride; // @[TensorUtil.scala 303:25:@6175.6]
  assign _GEN_34 = {{10'd0}, xfer_stride_pulses}; // @[TensorUtil.scala 305:16:@6178.8]
  assign _T_195 = xsize < _GEN_34; // @[TensorUtil.scala 305:16:@6178.8]
  assign _T_198 = xfer_stride_pulses - 9'h1; // @[TensorUtil.scala 309:33:@6184.10]
  assign _T_199 = $unsigned(_T_198); // @[TensorUtil.scala 309:33:@6185.10]
  assign _T_200 = _T_199[8:0]; // @[TensorUtil.scala 309:33:@6186.10]
  assign _T_201 = xsize - _GEN_34; // @[TensorUtil.scala 310:21:@6188.10]
  assign _T_202 = $unsigned(_T_201); // @[TensorUtil.scala 310:21:@6189.10]
  assign _T_203 = _T_202[18:0]; // @[TensorUtil.scala 310:21:@6190.10]
  assign _GEN_2 = _T_195 ? xsize : {{10'd0}, _T_200}; // @[TensorUtil.scala 305:38:@6179.8]
  assign _GEN_3 = _T_195 ? 19'h0 : _T_203; // @[TensorUtil.scala 305:38:@6179.8]
  assign _T_204 = io_xupdate & split; // @[TensorUtil.scala 312:25:@6195.8]
  assign _GEN_36 = {{7'd0}, xfer_split_pulses}; // @[TensorUtil.scala 314:15:@6198.10]
  assign _T_205 = xrem < _GEN_36; // @[TensorUtil.scala 314:15:@6198.10]
  assign _T_208 = xfer_split_pulses - 9'h1; // @[TensorUtil.scala 318:32:@6204.12]
  assign _T_209 = $unsigned(_T_208); // @[TensorUtil.scala 318:32:@6205.12]
  assign _T_210 = _T_209[8:0]; // @[TensorUtil.scala 318:32:@6206.12]
  assign _T_211 = xrem - _GEN_36; // @[TensorUtil.scala 319:20:@6208.12]
  assign _T_212 = $unsigned(_T_211); // @[TensorUtil.scala 319:20:@6209.12]
  assign _T_213 = _T_212[15:0]; // @[TensorUtil.scala 319:20:@6210.12]
  assign _GEN_4 = _T_205 ? xrem : {{7'd0}, _T_210}; // @[TensorUtil.scala 314:36:@6199.10]
  assign _GEN_5 = _T_205 ? 16'h0 : _T_213; // @[TensorUtil.scala 314:36:@6199.10]
  assign _GEN_6 = _T_204 ? {{20'd0}, xfer_split_bytes} : xfer_bytes; // @[TensorUtil.scala 312:35:@6196.8]
  assign _GEN_7 = _T_204 ? _GEN_4 : {{8'd0}, len}; // @[TensorUtil.scala 312:35:@6196.8]
  assign _GEN_8 = _T_204 ? _GEN_5 : xrem; // @[TensorUtil.scala 312:35:@6196.8]
  assign _GEN_9 = _T_194 ? {{20'd0}, xfer_stride_bytes} : _GEN_6; // @[TensorUtil.scala 303:36:@6176.6]
  assign _GEN_10 = _T_194 ? _GEN_2 : {{3'd0}, _GEN_7}; // @[TensorUtil.scala 303:36:@6176.6]
  assign _GEN_11 = _T_194 ? _GEN_3 : {{3'd0}, _GEN_8}; // @[TensorUtil.scala 303:36:@6176.6]
  assign _GEN_13 = io_start ? _GEN_0 : _GEN_10; // @[TensorUtil.scala 294:18:@6156.4]
  assign _GEN_14 = io_start ? _GEN_1 : _GEN_11; // @[TensorUtil.scala 294:18:@6156.4]
  assign _T_216 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@6219.8]
  assign _T_217 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@6220.8]
  assign _GEN_15 = io_xupdate ? _T_217 : xcnt; // @[TensorUtil.scala 325:26:@6218.6]
  assign _T_219 = io_yupdate & stride; // @[TensorUtil.scala 331:25:@6227.6]
  assign _T_221 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@6229.8]
  assign _T_222 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@6230.8]
  assign _GEN_17 = _T_219 ? _T_222 : ycnt; // @[TensorUtil.scala 331:36:@6228.6]
  assign _GEN_19 = stride ? xfer_stride_addr : caddr; // @[TensorUtil.scala 341:24:@6243.10]
  assign _GEN_20 = stride ? xfer_stride_addr : baddr; // @[TensorUtil.scala 341:24:@6243.10]
  assign _GEN_21 = split ? xfer_split_addr : _GEN_19; // @[TensorUtil.scala 339:17:@6239.8]
  assign _GEN_22 = split ? baddr : _GEN_20; // @[TensorUtil.scala 339:17:@6239.8]
  assign _GEN_23 = io_yupdate ? _GEN_21 : caddr; // @[TensorUtil.scala 338:26:@6238.6]
  assign _GEN_24 = io_yupdate ? _GEN_22 : baddr; // @[TensorUtil.scala 338:26:@6238.6]
  assign _GEN_25 = io_start ? xfer_init_addr : {{6'd0}, _GEN_23}; // @[TensorUtil.scala 335:18:@6233.4]
  assign _GEN_26 = io_start ? xfer_init_addr : {{6'd0}, _GEN_24}; // @[TensorUtil.scala 335:18:@6233.4]
  assign _T_232 = ycnt == _T_180; // @[TensorUtil.scala 354:10:@6260.4]
  assign io_done = _T_176 & _T_232; // @[TensorUtil.scala 352:11:@6262.4]
  assign io_stride = _T_176 & _T_181; // @[TensorUtil.scala 347:13:@6248.4]
  assign io_split = _T_173 & _T_184; // @[TensorUtil.scala 348:12:@6249.4]
  assign io_addr = caddr; // @[TensorUtil.scala 350:11:@6252.4]
  assign io_len = len; // @[TensorUtil.scala 351:10:@6253.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  caddr = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  baddr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  len = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  xcnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xrem = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ycnt = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  xfer_bytes = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    caddr <= _GEN_25[31:0];
    baddr <= _GEN_26[31:0];
    len <= _GEN_13[7:0];
    if (io_xinit) begin
      xcnt <= 8'h0;
    end else begin
      if (io_xupdate) begin
        xcnt <= _T_217;
      end
    end
    xrem <= _GEN_14[15:0];
    if (io_start) begin
      ycnt <= 16'h0;
    end else begin
      if (_T_219) begin
        ycnt <= _T_222;
      end
    end
    if (io_start) begin
      xfer_bytes <= {{20'd0}, xfer_init_bytes};
    end else begin
      if (_T_194) begin
        xfer_bytes <= {{20'd0}, xfer_stride_bytes};
      end else begin
        if (_T_204) begin
          xfer_bytes <= {{20'd0}, xfer_split_bytes};
        end
      end
    end
  end
endmodule
module TensorPadCtrl_8( // @[:@6264.2]
  input          clock, // @[:@6265.4]
  input          reset, // @[:@6266.4]
  input          io_start, // @[:@6267.4]
  output         io_done, // @[:@6267.4]
  input  [127:0] io_inst // @[:@6267.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@6292.4]
  wire [3:0] dec_ypad_0; // @[TensorUtil.scala 173:29:@6296.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@6300.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@6302.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@6304.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@6305.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@6306.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@6307.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@6308.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@6308.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@6309.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@6310.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@6310.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@6311.4]
  wire [18:0] _GEN_12; // @[TensorUtil.scala 182:46:@6312.4]
  wire [18:0] _T_39; // @[TensorUtil.scala 182:46:@6312.4]
  wire [19:0] _T_41; // @[TensorUtil.scala 182:71:@6313.4]
  wire [19:0] _T_42; // @[TensorUtil.scala 182:71:@6314.4]
  wire [18:0] xval; // @[TensorUtil.scala 182:71:@6315.4]
  wire  _T_44; // @[TensorUtil.scala 190:22:@6316.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 190:42:@6317.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 190:42:@6318.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 190:42:@6319.4]
  wire [3:0] yval; // @[TensorUtil.scala 190:10:@6320.4]
  reg  state; // @[TensorUtil.scala 197:22:@6321.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@6322.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@6324.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@6331.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@6332.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@6333.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@6334.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@6330.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@6323.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@6338.4]
  wire [18:0] _GEN_4; // @[TensorUtil.scala 212:25:@6339.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@6345.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@6352.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@6353.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@6351.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@6357.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@6358.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@6365.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@6367.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@6368.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@6366.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@6373.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@6292.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorUtil.scala 173:29:@6296.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@6300.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@6302.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@6308.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@6308.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@6309.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@6310.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@6310.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@6311.4]
  assign _GEN_12 = {{3'd0}, _T_38}; // @[TensorUtil.scala 182:46:@6312.4]
  assign _T_39 = _GEN_12 << 3; // @[TensorUtil.scala 182:46:@6312.4]
  assign _T_41 = _T_39 - 19'h1; // @[TensorUtil.scala 182:71:@6313.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@6314.4]
  assign xval = _T_42[18:0]; // @[TensorUtil.scala 182:71:@6315.4]
  assign _T_44 = dec_ypad_0 != 4'h0; // @[TensorUtil.scala 190:22:@6316.4]
  assign _T_46 = dec_ypad_0 - 4'h1; // @[TensorUtil.scala 190:42:@6317.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 190:42:@6318.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 190:42:@6319.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 190:10:@6320.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@6322.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@6324.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@6331.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@6332.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@6333.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@6334.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@6330.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@6323.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@6338.4]
  assign _GEN_4 = _T_56 ? xval : {{3'd0}, xmax}; // @[TensorUtil.scala 212:25:@6339.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@6345.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6352.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6353.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@6351.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@6357.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@6358.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@6365.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@6367.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@6368.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@6366.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@6373.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@6376.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_9( // @[:@6378.2]
  input          clock, // @[:@6379.4]
  input          reset, // @[:@6380.4]
  input          io_start, // @[:@6381.4]
  output         io_done, // @[:@6381.4]
  input  [127:0] io_inst // @[:@6381.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@6406.4]
  wire [3:0] dec_ypad_1; // @[TensorUtil.scala 173:29:@6412.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@6414.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@6416.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@6418.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@6419.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@6420.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@6421.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@6422.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@6422.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@6423.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@6424.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@6424.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@6425.4]
  wire [18:0] _GEN_12; // @[TensorUtil.scala 182:46:@6426.4]
  wire [18:0] _T_39; // @[TensorUtil.scala 182:46:@6426.4]
  wire [19:0] _T_41; // @[TensorUtil.scala 182:71:@6427.4]
  wire [19:0] _T_42; // @[TensorUtil.scala 182:71:@6428.4]
  wire [18:0] xval; // @[TensorUtil.scala 182:71:@6429.4]
  wire  _T_44; // @[TensorUtil.scala 192:22:@6430.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 192:42:@6431.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 192:42:@6432.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 192:42:@6433.4]
  wire [3:0] yval; // @[TensorUtil.scala 192:10:@6434.4]
  reg  state; // @[TensorUtil.scala 197:22:@6435.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@6436.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@6438.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@6445.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@6446.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@6447.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@6448.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@6444.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@6437.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@6452.4]
  wire [18:0] _GEN_4; // @[TensorUtil.scala 212:25:@6453.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@6459.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@6466.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@6467.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@6465.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@6471.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@6472.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@6479.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@6481.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@6482.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@6480.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@6487.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@6406.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorUtil.scala 173:29:@6412.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@6414.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@6416.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@6422.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@6422.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@6423.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@6424.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@6424.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@6425.4]
  assign _GEN_12 = {{3'd0}, _T_38}; // @[TensorUtil.scala 182:46:@6426.4]
  assign _T_39 = _GEN_12 << 3; // @[TensorUtil.scala 182:46:@6426.4]
  assign _T_41 = _T_39 - 19'h1; // @[TensorUtil.scala 182:71:@6427.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@6428.4]
  assign xval = _T_42[18:0]; // @[TensorUtil.scala 182:71:@6429.4]
  assign _T_44 = dec_ypad_1 != 4'h0; // @[TensorUtil.scala 192:22:@6430.4]
  assign _T_46 = dec_ypad_1 - 4'h1; // @[TensorUtil.scala 192:42:@6431.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 192:42:@6432.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 192:42:@6433.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 192:10:@6434.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@6436.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@6438.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@6445.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@6446.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@6447.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@6448.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@6444.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@6437.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@6452.4]
  assign _GEN_4 = _T_56 ? xval : {{3'd0}, xmax}; // @[TensorUtil.scala 212:25:@6453.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@6459.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6466.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6467.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@6465.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@6471.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@6472.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@6479.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@6481.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@6482.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@6480.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@6487.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@6490.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_10( // @[:@6492.2]
  input          clock, // @[:@6493.4]
  input          reset, // @[:@6494.4]
  input          io_start, // @[:@6495.4]
  output         io_done, // @[:@6495.4]
  input  [127:0] io_inst // @[:@6495.4]
);
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@6528.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@6532.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@6534.4]
  reg [31:0] _RAND_1;
  wire [6:0] _GEN_10; // @[TensorUtil.scala 184:19:@6536.4]
  wire [6:0] _T_35; // @[TensorUtil.scala 184:19:@6536.4]
  wire [7:0] _T_37; // @[TensorUtil.scala 184:44:@6537.4]
  wire [7:0] _T_38; // @[TensorUtil.scala 184:44:@6538.4]
  wire [6:0] xval; // @[TensorUtil.scala 184:44:@6539.4]
  reg  state; // @[TensorUtil.scala 197:22:@6540.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@6541.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@6543.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@6551.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@6553.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@6549.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@6542.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@6557.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@6564.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@6571.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@6572.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@6570.6]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@6528.4]
  assign _GEN_10 = {{3'd0}, dec_xpad_0}; // @[TensorUtil.scala 184:19:@6536.4]
  assign _T_35 = _GEN_10 << 3; // @[TensorUtil.scala 184:19:@6536.4]
  assign _T_37 = _T_35 - 7'h1; // @[TensorUtil.scala 184:44:@6537.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 184:44:@6538.4]
  assign xval = _T_38[6:0]; // @[TensorUtil.scala 184:44:@6539.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@6541.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@6543.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@6551.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@6553.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@6549.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@6542.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@6557.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@6564.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6571.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6572.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@6570.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@6595.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{9'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_11( // @[:@6597.2]
  input          clock, // @[:@6598.4]
  input          reset, // @[:@6599.4]
  input          io_start, // @[:@6600.4]
  output         io_done, // @[:@6600.4]
  input  [127:0] io_inst // @[:@6600.4]
);
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@6635.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@6637.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@6639.4]
  reg [31:0] _RAND_1;
  wire [6:0] _GEN_10; // @[TensorUtil.scala 186:19:@6641.4]
  wire [6:0] _T_35; // @[TensorUtil.scala 186:19:@6641.4]
  wire [7:0] _T_37; // @[TensorUtil.scala 186:44:@6642.4]
  wire [7:0] _T_38; // @[TensorUtil.scala 186:44:@6643.4]
  wire [6:0] xval; // @[TensorUtil.scala 186:44:@6644.4]
  reg  state; // @[TensorUtil.scala 197:22:@6645.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@6646.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@6648.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@6656.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@6658.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@6654.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@6647.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@6662.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@6669.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@6676.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@6677.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@6675.6]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@6635.4]
  assign _GEN_10 = {{3'd0}, dec_xpad_1}; // @[TensorUtil.scala 186:19:@6641.4]
  assign _T_35 = _GEN_10 << 3; // @[TensorUtil.scala 186:19:@6641.4]
  assign _T_37 = _T_35 - 7'h1; // @[TensorUtil.scala 186:44:@6642.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 186:44:@6643.4]
  assign xval = _T_38[6:0]; // @[TensorUtil.scala 186:44:@6644.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@6646.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@6648.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@6656.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@6658.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@6654.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@6647.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@6662.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@6669.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6676.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6677.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@6675.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@6700.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{9'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorLoad_2( // @[:@6702.2]
  input          clock, // @[:@6703.4]
  input          reset, // @[:@6704.4]
  input          io_start, // @[:@6705.4]
  output         io_done, // @[:@6705.4]
  input  [127:0] io_inst, // @[:@6705.4]
  input  [31:0]  io_baddr, // @[:@6705.4]
  input          io_vme_rd_cmd_ready, // @[:@6705.4]
  output         io_vme_rd_cmd_valid, // @[:@6705.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@6705.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@6705.4]
  output         io_vme_rd_data_ready, // @[:@6705.4]
  input          io_vme_rd_data_valid, // @[:@6705.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@6705.4]
  input          io_tensor_rd_idx_valid, // @[:@6705.4]
  input  [10:0]  io_tensor_rd_idx_bits, // @[:@6705.4]
  output         io_tensor_rd_data_valid, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_0, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_1, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_2, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_3, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_4, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_5, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_6, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_7, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_8, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_9, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_10, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_11, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_12, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_13, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_14, // @[:@6705.4]
  output [31:0]  io_tensor_rd_data_bits_0_15, // @[:@6705.4]
  input          io_tensor_wr_valid, // @[:@6705.4]
  input  [10:0]  io_tensor_wr_bits_idx, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_0, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_1, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_2, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_3, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_4, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_5, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_6, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_7, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_8, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_9, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_10, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_11, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_12, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_13, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_14, // @[:@6705.4]
  input  [31:0]  io_tensor_wr_bits_data_0_15 // @[:@6705.4]
);
  wire  dataCtrl_clock; // @[TensorLoad.scala 52:24:@6742.4]
  wire  dataCtrl_io_start; // @[TensorLoad.scala 52:24:@6742.4]
  wire  dataCtrl_io_done; // @[TensorLoad.scala 52:24:@6742.4]
  wire [127:0] dataCtrl_io_inst; // @[TensorLoad.scala 52:24:@6742.4]
  wire [31:0] dataCtrl_io_baddr; // @[TensorLoad.scala 52:24:@6742.4]
  wire  dataCtrl_io_xinit; // @[TensorLoad.scala 52:24:@6742.4]
  wire  dataCtrl_io_xupdate; // @[TensorLoad.scala 52:24:@6742.4]
  wire  dataCtrl_io_yupdate; // @[TensorLoad.scala 52:24:@6742.4]
  wire  dataCtrl_io_stride; // @[TensorLoad.scala 52:24:@6742.4]
  wire  dataCtrl_io_split; // @[TensorLoad.scala 52:24:@6742.4]
  wire [31:0] dataCtrl_io_addr; // @[TensorLoad.scala 52:24:@6742.4]
  wire [7:0] dataCtrl_io_len; // @[TensorLoad.scala 52:24:@6742.4]
  wire  yPadCtrl0_clock; // @[TensorLoad.scala 55:25:@6746.4]
  wire  yPadCtrl0_reset; // @[TensorLoad.scala 55:25:@6746.4]
  wire  yPadCtrl0_io_start; // @[TensorLoad.scala 55:25:@6746.4]
  wire  yPadCtrl0_io_done; // @[TensorLoad.scala 55:25:@6746.4]
  wire [127:0] yPadCtrl0_io_inst; // @[TensorLoad.scala 55:25:@6746.4]
  wire  yPadCtrl1_clock; // @[TensorLoad.scala 56:25:@6749.4]
  wire  yPadCtrl1_reset; // @[TensorLoad.scala 56:25:@6749.4]
  wire  yPadCtrl1_io_start; // @[TensorLoad.scala 56:25:@6749.4]
  wire  yPadCtrl1_io_done; // @[TensorLoad.scala 56:25:@6749.4]
  wire [127:0] yPadCtrl1_io_inst; // @[TensorLoad.scala 56:25:@6749.4]
  wire  xPadCtrl0_clock; // @[TensorLoad.scala 57:25:@6752.4]
  wire  xPadCtrl0_reset; // @[TensorLoad.scala 57:25:@6752.4]
  wire  xPadCtrl0_io_start; // @[TensorLoad.scala 57:25:@6752.4]
  wire  xPadCtrl0_io_done; // @[TensorLoad.scala 57:25:@6752.4]
  wire [127:0] xPadCtrl0_io_inst; // @[TensorLoad.scala 57:25:@6752.4]
  wire  xPadCtrl1_clock; // @[TensorLoad.scala 58:25:@6755.4]
  wire  xPadCtrl1_reset; // @[TensorLoad.scala 58:25:@6755.4]
  wire  xPadCtrl1_io_start; // @[TensorLoad.scala 58:25:@6755.4]
  wire  xPadCtrl1_io_done; // @[TensorLoad.scala 58:25:@6755.4]
  wire [127:0] xPadCtrl1_io_inst; // @[TensorLoad.scala 58:25:@6755.4]
  reg [63:0] tensorFile_0_0 [0:2047]; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] _RAND_0;
  wire [63:0] tensorFile_0_0_rdata_0_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_0_rdata_0_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire [63:0] tensorFile_0_0__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_0__T_992_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_0__T_992_mask; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_0__T_992_en; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] tensorFile_0_1 [0:2047]; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] _RAND_1;
  wire [63:0] tensorFile_0_1_rdata_0_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_1_rdata_0_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire [63:0] tensorFile_0_1__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_1__T_992_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_1__T_992_mask; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_1__T_992_en; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] tensorFile_0_2 [0:2047]; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] _RAND_2;
  wire [63:0] tensorFile_0_2_rdata_0_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_2_rdata_0_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire [63:0] tensorFile_0_2__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_2__T_992_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_2__T_992_mask; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_2__T_992_en; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] tensorFile_0_3 [0:2047]; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] _RAND_3;
  wire [63:0] tensorFile_0_3_rdata_0_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_3_rdata_0_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire [63:0] tensorFile_0_3__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_3__T_992_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_3__T_992_mask; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_3__T_992_en; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] tensorFile_0_4 [0:2047]; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] _RAND_4;
  wire [63:0] tensorFile_0_4_rdata_0_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_4_rdata_0_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire [63:0] tensorFile_0_4__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_4__T_992_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_4__T_992_mask; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_4__T_992_en; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] tensorFile_0_5 [0:2047]; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] _RAND_5;
  wire [63:0] tensorFile_0_5_rdata_0_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_5_rdata_0_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire [63:0] tensorFile_0_5__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_5__T_992_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_5__T_992_mask; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_5__T_992_en; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] tensorFile_0_6 [0:2047]; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] _RAND_6;
  wire [63:0] tensorFile_0_6_rdata_0_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_6_rdata_0_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire [63:0] tensorFile_0_6__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_6__T_992_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_6__T_992_mask; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_6__T_992_en; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] tensorFile_0_7 [0:2047]; // @[TensorLoad.scala 222:16:@7025.4]
  reg [63:0] _RAND_7;
  wire [63:0] tensorFile_0_7_rdata_0_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_7_rdata_0_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire [63:0] tensorFile_0_7__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
  wire [10:0] tensorFile_0_7__T_992_addr; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_7__T_992_mask; // @[TensorLoad.scala 222:16:@7025.4]
  wire  tensorFile_0_7__T_992_en; // @[TensorLoad.scala 222:16:@7025.4]
  wire [15:0] dec_sram_offset; // @[TensorLoad.scala 51:29:@6722.4]
  wire [15:0] dec_xsize; // @[TensorLoad.scala 51:29:@6730.4]
  wire [3:0] dec_ypad_0; // @[TensorLoad.scala 51:29:@6734.4]
  wire [3:0] dec_ypad_1; // @[TensorLoad.scala 51:29:@6736.4]
  wire [3:0] dec_xpad_0; // @[TensorLoad.scala 51:29:@6738.4]
  wire [3:0] dec_xpad_1; // @[TensorLoad.scala 51:29:@6740.4]
  reg  dataCtrlDone; // @[TensorLoad.scala 54:29:@6745.4]
  reg [31:0] _RAND_8;
  reg [2:0] tag; // @[TensorLoad.scala 60:16:@6758.4]
  reg [31:0] _RAND_9;
  reg [2:0] state; // @[TensorLoad.scala 65:22:@6760.4]
  reg [31:0] _RAND_10;
  wire  _T_614; // @[Conditional.scala 37:30:@6761.4]
  wire  _T_616; // @[TensorLoad.scala 71:25:@6764.8]
  wire  _T_618; // @[TensorLoad.scala 73:31:@6769.10]
  wire [2:0] _GEN_0; // @[TensorLoad.scala 73:40:@6770.10]
  wire [2:0] _GEN_1; // @[TensorLoad.scala 71:34:@6765.8]
  wire [2:0] _GEN_2; // @[TensorLoad.scala 70:22:@6763.6]
  wire  _T_619; // @[Conditional.scala 37:30:@6779.6]
  wire [2:0] _GEN_4; // @[TensorLoad.scala 81:31:@6781.8]
  wire  _T_622; // @[Conditional.scala 37:30:@6792.8]
  wire [2:0] _GEN_5; // @[TensorLoad.scala 90:31:@6794.10]
  wire  _T_623; // @[Conditional.scala 37:30:@6799.10]
  wire [2:0] _GEN_6; // @[TensorLoad.scala 95:33:@6801.12]
  wire  _T_624; // @[Conditional.scala 37:30:@6806.12]
  wire  _T_626; // @[TensorLoad.scala 102:27:@6810.18]
  wire  _T_628; // @[TensorLoad.scala 104:33:@6815.20]
  wire [2:0] _GEN_7; // @[TensorLoad.scala 104:42:@6816.20]
  wire [2:0] _GEN_8; // @[TensorLoad.scala 102:36:@6811.18]
  wire [2:0] _GEN_10; // @[TensorLoad.scala 110:36:@6826.20]
  wire [2:0] _GEN_11; // @[TensorLoad.scala 117:39:@6839.20]
  wire [2:0] _GEN_12; // @[TensorLoad.scala 109:40:@6824.18]
  wire [2:0] _GEN_13; // @[TensorLoad.scala 101:32:@6809.16]
  wire [2:0] _GEN_14; // @[TensorLoad.scala 100:34:@6808.14]
  wire  _T_633; // @[Conditional.scala 37:30:@6845.14]
  wire [2:0] _GEN_17; // @[TensorLoad.scala 124:28:@6848.18]
  wire [2:0] _GEN_18; // @[TensorLoad.scala 123:31:@6847.16]
  wire  _T_638; // @[Conditional.scala 37:30:@6869.16]
  wire  _T_639; // @[TensorLoad.scala 140:30:@6871.18]
  wire [2:0] _GEN_19; // @[TensorLoad.scala 140:47:@6872.18]
  wire [2:0] _GEN_20; // @[Conditional.scala 39:67:@6870.16]
  wire [2:0] _GEN_21; // @[Conditional.scala 39:67:@6846.14]
  wire [2:0] _GEN_22; // @[Conditional.scala 39:67:@6807.12]
  wire [2:0] _GEN_23; // @[Conditional.scala 39:67:@6800.10]
  wire [2:0] _GEN_24; // @[Conditional.scala 39:67:@6793.8]
  wire [2:0] _GEN_25; // @[Conditional.scala 39:67:@6780.6]
  wire [2:0] _GEN_26; // @[Conditional.scala 40:58:@6762.4]
  wire  _T_640; // @[TensorLoad.scala 147:30:@6876.4]
  wire  _T_641; // @[TensorLoad.scala 147:40:@6877.4]
  wire  _T_643; // @[Decoupled.scala 37:37:@6883.4]
  wire  _T_648; // @[TensorLoad.scala 156:36:@6893.6]
  wire  _GEN_27; // @[TensorLoad.scala 156:57:@6894.6]
  wire  _GEN_28; // @[TensorLoad.scala 154:25:@6888.4]
  wire  _T_653; // @[TensorLoad.scala 161:44:@6899.4]
  wire  _T_660; // @[TensorLoad.scala 164:61:@6905.4]
  wire  _T_661; // @[TensorLoad.scala 164:48:@6906.4]
  wire  _T_662; // @[TensorLoad.scala 165:14:@6907.4]
  wire  _T_663; // @[TensorLoad.scala 165:25:@6908.4]
  wire  _T_664; // @[TensorLoad.scala 165:45:@6909.4]
  wire  _T_665; // @[TensorLoad.scala 164:70:@6910.4]
  wire  _T_671; // @[TensorLoad.scala 169:14:@6916.4]
  wire  _T_672; // @[TensorLoad.scala 169:25:@6917.4]
  wire  _T_673; // @[TensorLoad.scala 168:35:@6918.4]
  wire  _T_675; // @[TensorLoad.scala 170:32:@6920.4]
  wire  _T_676; // @[TensorLoad.scala 170:30:@6921.4]
  wire  _T_677; // @[TensorLoad.scala 170:46:@6922.4]
  wire  _T_680; // @[TensorLoad.scala 170:67:@6924.4]
  wire  _T_681; // @[TensorLoad.scala 169:46:@6925.4]
  wire  _T_685; // @[TensorLoad.scala 171:45:@6929.4]
  wire  _T_686; // @[TensorLoad.scala 170:89:@6930.4]
  wire  _T_691; // @[TensorLoad.scala 173:44:@6935.4]
  wire  _T_692; // @[TensorLoad.scala 174:28:@6936.4]
  wire  _T_693; // @[TensorLoad.scala 174:46:@6937.4]
  wire  _T_696; // @[TensorLoad.scala 174:67:@6939.4]
  wire  _T_697; // @[TensorLoad.scala 174:25:@6940.4]
  wire  _T_699; // @[TensorLoad.scala 182:32:@6947.4]
  wire  _T_702; // @[TensorLoad.scala 190:11:@6954.4]
  wire  _T_703; // @[TensorLoad.scala 189:36:@6955.4]
  wire  _T_705; // @[TensorLoad.scala 190:22:@6957.4]
  wire  _T_706; // @[TensorLoad.scala 192:11:@6958.4]
  wire  isZeroPad; // @[TensorLoad.scala 191:22:@6959.4]
  wire  _T_709; // @[TensorLoad.scala 194:24:@6962.4]
  wire  _T_711; // @[TensorLoad.scala 194:53:@6963.4]
  wire  _T_712; // @[TensorLoad.scala 194:46:@6964.4]
  wire  _T_715; // @[TensorLoad.scala 196:36:@6970.6]
  wire [3:0] _T_717; // @[TensorLoad.scala 197:16:@6972.8]
  wire [2:0] _T_718; // @[TensorLoad.scala 197:16:@6973.8]
  wire [2:0] _GEN_29; // @[TensorLoad.scala 196:50:@6971.6]
  wire  _T_732; // @[TensorLoad.scala 202:51:@6989.6]
  reg [10:0] waddr_cur; // @[TensorLoad.scala 206:22:@6995.4]
  reg [31:0] _RAND_11;
  reg [10:0] waddr_nxt; // @[TensorLoad.scala 207:22:@6996.4]
  reg [31:0] _RAND_12;
  wire [11:0] _T_748; // @[TensorLoad.scala 215:28:@7010.8]
  wire [10:0] _T_749; // @[TensorLoad.scala 215:28:@7011.8]
  wire  _T_751; // @[TensorLoad.scala 216:33:@7016.8]
  wire [15:0] _GEN_126; // @[TensorLoad.scala 217:28:@7018.10]
  wire [16:0] _T_752; // @[TensorLoad.scala 217:28:@7018.10]
  wire [15:0] _T_753; // @[TensorLoad.scala 217:28:@7019.10]
  wire [15:0] _GEN_33; // @[TensorLoad.scala 216:59:@7017.8]
  wire [15:0] _GEN_34; // @[TensorLoad.scala 216:59:@7017.8]
  wire [15:0] _GEN_35; // @[TensorLoad.scala 214:3:@7009.6]
  wire [15:0] _GEN_36; // @[TensorLoad.scala 214:3:@7009.6]
  wire [15:0] _GEN_37; // @[TensorLoad.scala 208:25:@6998.4]
  wire [15:0] _GEN_38; // @[TensorLoad.scala 208:25:@6998.4]
  wire  wmask_0_0; // @[TensorLoad.scala 235:26:@7037.4]
  wire [63:0] wdata_0_0; // @[TensorLoad.scala 236:25:@7039.4]
  wire  wmask_0_1; // @[TensorLoad.scala 235:26:@7041.4]
  wire  wmask_0_2; // @[TensorLoad.scala 235:26:@7045.4]
  wire  wmask_0_3; // @[TensorLoad.scala 235:26:@7049.4]
  wire  wmask_0_4; // @[TensorLoad.scala 235:26:@7053.4]
  wire  wmask_0_5; // @[TensorLoad.scala 235:26:@7057.4]
  wire  wmask_0_6; // @[TensorLoad.scala 235:26:@7061.4]
  wire [255:0] _T_855; // @[TensorLoad.scala 238:43:@7075.4]
  wire [511:0] _T_863; // @[TensorLoad.scala 238:43:@7083.4]
  wire [63:0] _T_915; // @[TensorLoad.scala 238:58:@7087.4]
  wire [63:0] _T_916; // @[TensorLoad.scala 238:58:@7089.4]
  wire [63:0] _T_917; // @[TensorLoad.scala 238:58:@7091.4]
  wire [63:0] _T_918; // @[TensorLoad.scala 238:58:@7093.4]
  wire [63:0] _T_919; // @[TensorLoad.scala 238:58:@7095.4]
  wire [63:0] _T_920; // @[TensorLoad.scala 238:58:@7097.4]
  wire [63:0] _T_921; // @[TensorLoad.scala 238:58:@7099.4]
  wire [63:0] _T_922; // @[TensorLoad.scala 238:58:@7101.4]
  reg  rvalid; // @[TensorLoad.scala 252:23:@7142.4]
  reg [31:0] _RAND_13;
  wire  _GEN_75; // @[TensorLoad.scala 256:26:@7147.4]
  wire [511:0] _T_1043; // @[TensorLoad.scala 259:38:@7159.4]
  wire  _T_1191; // @[TensorLoad.scala 263:96:@7215.4]
  wire  done_no_pad; // @[TensorLoad.scala 263:83:@7216.4]
  wire  done_x_pad; // @[TensorLoad.scala 264:72:@7221.4]
  wire  _T_1198; // @[TensorLoad.scala 265:37:@7223.4]
  wire  done_y_pad; // @[TensorLoad.scala 265:52:@7224.4]
  wire  _T_1199; // @[TensorLoad.scala 266:26:@7225.4]
  reg [10:0] tensorFile_0_0_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [10:0] tensorFile_0_1_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [10:0] tensorFile_0_2_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_16;
  reg [10:0] tensorFile_0_3_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [10:0] tensorFile_0_4_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_18;
  reg [10:0] tensorFile_0_5_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [10:0] tensorFile_0_6_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_20;
  reg [10:0] tensorFile_0_7_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_21;
  TensorDataCtrl_2 dataCtrl ( // @[TensorLoad.scala 52:24:@6742.4]
    .clock(dataCtrl_clock),
    .io_start(dataCtrl_io_start),
    .io_done(dataCtrl_io_done),
    .io_inst(dataCtrl_io_inst),
    .io_baddr(dataCtrl_io_baddr),
    .io_xinit(dataCtrl_io_xinit),
    .io_xupdate(dataCtrl_io_xupdate),
    .io_yupdate(dataCtrl_io_yupdate),
    .io_stride(dataCtrl_io_stride),
    .io_split(dataCtrl_io_split),
    .io_addr(dataCtrl_io_addr),
    .io_len(dataCtrl_io_len)
  );
  TensorPadCtrl_8 yPadCtrl0 ( // @[TensorLoad.scala 55:25:@6746.4]
    .clock(yPadCtrl0_clock),
    .reset(yPadCtrl0_reset),
    .io_start(yPadCtrl0_io_start),
    .io_done(yPadCtrl0_io_done),
    .io_inst(yPadCtrl0_io_inst)
  );
  TensorPadCtrl_9 yPadCtrl1 ( // @[TensorLoad.scala 56:25:@6749.4]
    .clock(yPadCtrl1_clock),
    .reset(yPadCtrl1_reset),
    .io_start(yPadCtrl1_io_start),
    .io_done(yPadCtrl1_io_done),
    .io_inst(yPadCtrl1_io_inst)
  );
  TensorPadCtrl_10 xPadCtrl0 ( // @[TensorLoad.scala 57:25:@6752.4]
    .clock(xPadCtrl0_clock),
    .reset(xPadCtrl0_reset),
    .io_start(xPadCtrl0_io_start),
    .io_done(xPadCtrl0_io_done),
    .io_inst(xPadCtrl0_io_inst)
  );
  TensorPadCtrl_11 xPadCtrl1 ( // @[TensorLoad.scala 58:25:@6755.4]
    .clock(xPadCtrl1_clock),
    .reset(xPadCtrl1_reset),
    .io_start(xPadCtrl1_io_start),
    .io_done(xPadCtrl1_io_done),
    .io_inst(xPadCtrl1_io_inst)
  );
  assign tensorFile_0_0_rdata_0_addr = tensorFile_0_0_rdata_0_addr_pipe_0;
  assign tensorFile_0_0_rdata_0_data = tensorFile_0_0[tensorFile_0_0_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7025.4]
  assign tensorFile_0_0__T_992_data = _T_640 ? _T_915 : wdata_0_0;
  assign tensorFile_0_0__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_0__T_992_mask = _T_640 ? 1'h1 : wmask_0_0;
  assign tensorFile_0_0__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_1_rdata_0_addr = tensorFile_0_1_rdata_0_addr_pipe_0;
  assign tensorFile_0_1_rdata_0_data = tensorFile_0_1[tensorFile_0_1_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7025.4]
  assign tensorFile_0_1__T_992_data = _T_640 ? _T_916 : wdata_0_0;
  assign tensorFile_0_1__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_1__T_992_mask = _T_640 ? 1'h1 : wmask_0_1;
  assign tensorFile_0_1__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_2_rdata_0_addr = tensorFile_0_2_rdata_0_addr_pipe_0;
  assign tensorFile_0_2_rdata_0_data = tensorFile_0_2[tensorFile_0_2_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7025.4]
  assign tensorFile_0_2__T_992_data = _T_640 ? _T_917 : wdata_0_0;
  assign tensorFile_0_2__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_2__T_992_mask = _T_640 ? 1'h1 : wmask_0_2;
  assign tensorFile_0_2__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_3_rdata_0_addr = tensorFile_0_3_rdata_0_addr_pipe_0;
  assign tensorFile_0_3_rdata_0_data = tensorFile_0_3[tensorFile_0_3_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7025.4]
  assign tensorFile_0_3__T_992_data = _T_640 ? _T_918 : wdata_0_0;
  assign tensorFile_0_3__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_3__T_992_mask = _T_640 ? 1'h1 : wmask_0_3;
  assign tensorFile_0_3__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_4_rdata_0_addr = tensorFile_0_4_rdata_0_addr_pipe_0;
  assign tensorFile_0_4_rdata_0_data = tensorFile_0_4[tensorFile_0_4_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7025.4]
  assign tensorFile_0_4__T_992_data = _T_640 ? _T_919 : wdata_0_0;
  assign tensorFile_0_4__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_4__T_992_mask = _T_640 ? 1'h1 : wmask_0_4;
  assign tensorFile_0_4__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_5_rdata_0_addr = tensorFile_0_5_rdata_0_addr_pipe_0;
  assign tensorFile_0_5_rdata_0_data = tensorFile_0_5[tensorFile_0_5_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7025.4]
  assign tensorFile_0_5__T_992_data = _T_640 ? _T_920 : wdata_0_0;
  assign tensorFile_0_5__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_5__T_992_mask = _T_640 ? 1'h1 : wmask_0_5;
  assign tensorFile_0_5__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_6_rdata_0_addr = tensorFile_0_6_rdata_0_addr_pipe_0;
  assign tensorFile_0_6_rdata_0_data = tensorFile_0_6[tensorFile_0_6_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7025.4]
  assign tensorFile_0_6__T_992_data = _T_640 ? _T_921 : wdata_0_0;
  assign tensorFile_0_6__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_6__T_992_mask = _T_640 ? 1'h1 : wmask_0_6;
  assign tensorFile_0_6__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_7_rdata_0_addr = tensorFile_0_7_rdata_0_addr_pipe_0;
  assign tensorFile_0_7_rdata_0_data = tensorFile_0_7[tensorFile_0_7_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7025.4]
  assign tensorFile_0_7__T_992_data = _T_640 ? _T_922 : wdata_0_0;
  assign tensorFile_0_7__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_7__T_992_mask = _T_640 ? 1'h1 : _T_711;
  assign tensorFile_0_7__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign dec_sram_offset = io_inst[24:9]; // @[TensorLoad.scala 51:29:@6722.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorLoad.scala 51:29:@6730.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorLoad.scala 51:29:@6734.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorLoad.scala 51:29:@6736.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorLoad.scala 51:29:@6738.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorLoad.scala 51:29:@6740.4]
  assign _T_614 = 3'h0 == state; // @[Conditional.scala 37:30:@6761.4]
  assign _T_616 = dec_ypad_0 != 4'h0; // @[TensorLoad.scala 71:25:@6764.8]
  assign _T_618 = dec_xpad_0 != 4'h0; // @[TensorLoad.scala 73:31:@6769.10]
  assign _GEN_0 = _T_618 ? 3'h2 : 3'h3; // @[TensorLoad.scala 73:40:@6770.10]
  assign _GEN_1 = _T_616 ? 3'h1 : _GEN_0; // @[TensorLoad.scala 71:34:@6765.8]
  assign _GEN_2 = io_start ? _GEN_1 : state; // @[TensorLoad.scala 70:22:@6763.6]
  assign _T_619 = 3'h1 == state; // @[Conditional.scala 37:30:@6779.6]
  assign _GEN_4 = yPadCtrl0_io_done ? _GEN_0 : state; // @[TensorLoad.scala 81:31:@6781.8]
  assign _T_622 = 3'h2 == state; // @[Conditional.scala 37:30:@6792.8]
  assign _GEN_5 = xPadCtrl0_io_done ? 3'h3 : state; // @[TensorLoad.scala 90:31:@6794.10]
  assign _T_623 = 3'h3 == state; // @[Conditional.scala 37:30:@6799.10]
  assign _GEN_6 = io_vme_rd_cmd_ready ? 3'h4 : state; // @[TensorLoad.scala 95:33:@6801.12]
  assign _T_624 = 3'h4 == state; // @[Conditional.scala 37:30:@6806.12]
  assign _T_626 = dec_xpad_1 != 4'h0; // @[TensorLoad.scala 102:27:@6810.18]
  assign _T_628 = dec_ypad_1 != 4'h0; // @[TensorLoad.scala 104:33:@6815.20]
  assign _GEN_7 = _T_628 ? 3'h6 : 3'h0; // @[TensorLoad.scala 104:42:@6816.20]
  assign _GEN_8 = _T_626 ? 3'h5 : _GEN_7; // @[TensorLoad.scala 102:36:@6811.18]
  assign _GEN_10 = _T_626 ? 3'h5 : _GEN_0; // @[TensorLoad.scala 110:36:@6826.20]
  assign _GEN_11 = dataCtrl_io_split ? 3'h3 : state; // @[TensorLoad.scala 117:39:@6839.20]
  assign _GEN_12 = dataCtrl_io_stride ? _GEN_10 : _GEN_11; // @[TensorLoad.scala 109:40:@6824.18]
  assign _GEN_13 = dataCtrl_io_done ? _GEN_8 : _GEN_12; // @[TensorLoad.scala 101:32:@6809.16]
  assign _GEN_14 = io_vme_rd_data_valid ? _GEN_13 : state; // @[TensorLoad.scala 100:34:@6808.14]
  assign _T_633 = 3'h5 == state; // @[Conditional.scala 37:30:@6845.14]
  assign _GEN_17 = dataCtrlDone ? _GEN_7 : _GEN_0; // @[TensorLoad.scala 124:28:@6848.18]
  assign _GEN_18 = xPadCtrl1_io_done ? _GEN_17 : state; // @[TensorLoad.scala 123:31:@6847.16]
  assign _T_638 = 3'h6 == state; // @[Conditional.scala 37:30:@6869.16]
  assign _T_639 = yPadCtrl1_io_done & dataCtrlDone; // @[TensorLoad.scala 140:30:@6871.18]
  assign _GEN_19 = _T_639 ? 3'h0 : state; // @[TensorLoad.scala 140:47:@6872.18]
  assign _GEN_20 = _T_638 ? _GEN_19 : state; // @[Conditional.scala 39:67:@6870.16]
  assign _GEN_21 = _T_633 ? _GEN_18 : _GEN_20; // @[Conditional.scala 39:67:@6846.14]
  assign _GEN_22 = _T_624 ? _GEN_14 : _GEN_21; // @[Conditional.scala 39:67:@6807.12]
  assign _GEN_23 = _T_623 ? _GEN_6 : _GEN_22; // @[Conditional.scala 39:67:@6800.10]
  assign _GEN_24 = _T_622 ? _GEN_5 : _GEN_23; // @[Conditional.scala 39:67:@6793.8]
  assign _GEN_25 = _T_619 ? _GEN_4 : _GEN_24; // @[Conditional.scala 39:67:@6780.6]
  assign _GEN_26 = _T_614 ? _GEN_2 : _GEN_25; // @[Conditional.scala 40:58:@6762.4]
  assign _T_640 = state == 3'h0; // @[TensorLoad.scala 147:30:@6876.4]
  assign _T_641 = _T_640 & io_start; // @[TensorLoad.scala 147:40:@6877.4]
  assign _T_643 = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[Decoupled.scala 37:37:@6883.4]
  assign _T_648 = _T_643 & dataCtrl_io_done; // @[TensorLoad.scala 156:36:@6893.6]
  assign _GEN_27 = _T_648 ? 1'h1 : dataCtrlDone; // @[TensorLoad.scala 156:57:@6894.6]
  assign _GEN_28 = _T_640 ? 1'h0 : _GEN_27; // @[TensorLoad.scala 154:25:@6888.4]
  assign _T_653 = _T_616 & _T_640; // @[TensorLoad.scala 161:44:@6899.4]
  assign _T_660 = dec_xpad_1 == 4'h0; // @[TensorLoad.scala 164:61:@6905.4]
  assign _T_661 = _T_648 & _T_660; // @[TensorLoad.scala 164:48:@6906.4]
  assign _T_662 = state == 3'h5; // @[TensorLoad.scala 165:14:@6907.4]
  assign _T_663 = _T_662 & xPadCtrl1_io_done; // @[TensorLoad.scala 165:25:@6908.4]
  assign _T_664 = _T_663 & dataCtrlDone; // @[TensorLoad.scala 165:45:@6909.4]
  assign _T_665 = _T_661 | _T_664; // @[TensorLoad.scala 164:70:@6910.4]
  assign _T_671 = state == 3'h1; // @[TensorLoad.scala 169:14:@6916.4]
  assign _T_672 = _T_671 & yPadCtrl0_io_done; // @[TensorLoad.scala 169:25:@6917.4]
  assign _T_673 = _T_641 | _T_672; // @[TensorLoad.scala 168:35:@6918.4]
  assign _T_675 = ~ dataCtrlDone; // @[TensorLoad.scala 170:32:@6920.4]
  assign _T_676 = _T_643 & _T_675; // @[TensorLoad.scala 170:30:@6921.4]
  assign _T_677 = _T_676 & dataCtrl_io_stride; // @[TensorLoad.scala 170:46:@6922.4]
  assign _T_680 = _T_677 & _T_660; // @[TensorLoad.scala 170:67:@6924.4]
  assign _T_681 = _T_673 | _T_680; // @[TensorLoad.scala 169:46:@6925.4]
  assign _T_685 = _T_663 & _T_675; // @[TensorLoad.scala 171:45:@6929.4]
  assign _T_686 = _T_681 | _T_685; // @[TensorLoad.scala 170:89:@6930.4]
  assign _T_691 = _T_626 & _T_643; // @[TensorLoad.scala 173:44:@6935.4]
  assign _T_692 = ~ dataCtrl_io_done; // @[TensorLoad.scala 174:28:@6936.4]
  assign _T_693 = _T_692 & dataCtrl_io_stride; // @[TensorLoad.scala 174:46:@6937.4]
  assign _T_696 = _T_693 & _T_626; // @[TensorLoad.scala 174:67:@6939.4]
  assign _T_697 = dataCtrl_io_done | _T_696; // @[TensorLoad.scala 174:25:@6940.4]
  assign _T_699 = state == 3'h3; // @[TensorLoad.scala 182:32:@6947.4]
  assign _T_702 = state == 3'h2; // @[TensorLoad.scala 190:11:@6954.4]
  assign _T_703 = _T_671 | _T_702; // @[TensorLoad.scala 189:36:@6955.4]
  assign _T_705 = _T_703 | _T_662; // @[TensorLoad.scala 190:22:@6957.4]
  assign _T_706 = state == 3'h6; // @[TensorLoad.scala 192:11:@6958.4]
  assign isZeroPad = _T_705 | _T_706; // @[TensorLoad.scala 191:22:@6959.4]
  assign _T_709 = _T_640 | _T_699; // @[TensorLoad.scala 194:24:@6962.4]
  assign _T_711 = tag == 3'h7; // @[TensorLoad.scala 194:53:@6963.4]
  assign _T_712 = _T_709 | _T_711; // @[TensorLoad.scala 194:46:@6964.4]
  assign _T_715 = _T_643 | isZeroPad; // @[TensorLoad.scala 196:36:@6970.6]
  assign _T_717 = tag + 3'h1; // @[TensorLoad.scala 197:16:@6972.8]
  assign _T_718 = tag + 3'h1; // @[TensorLoad.scala 197:16:@6973.8]
  assign _GEN_29 = _T_715 ? _T_718 : tag; // @[TensorLoad.scala 196:50:@6971.6]
  assign _T_732 = _T_715 & _T_711; // @[TensorLoad.scala 202:51:@6989.6]
  assign _T_748 = waddr_cur + 11'h1; // @[TensorLoad.scala 215:28:@7010.8]
  assign _T_749 = waddr_cur + 11'h1; // @[TensorLoad.scala 215:28:@7011.8]
  assign _T_751 = dataCtrl_io_stride & _T_643; // @[TensorLoad.scala 216:33:@7016.8]
  assign _GEN_126 = {{5'd0}, waddr_nxt}; // @[TensorLoad.scala 217:28:@7018.10]
  assign _T_752 = _GEN_126 + dec_xsize; // @[TensorLoad.scala 217:28:@7018.10]
  assign _T_753 = _GEN_126 + dec_xsize; // @[TensorLoad.scala 217:28:@7019.10]
  assign _GEN_33 = _T_751 ? _T_753 : {{5'd0}, waddr_cur}; // @[TensorLoad.scala 216:59:@7017.8]
  assign _GEN_34 = _T_751 ? _T_753 : {{5'd0}, waddr_nxt}; // @[TensorLoad.scala 216:59:@7017.8]
  assign _GEN_35 = _T_732 ? {{5'd0}, _T_749} : _GEN_33; // @[TensorLoad.scala 214:3:@7009.6]
  assign _GEN_36 = _T_732 ? {{5'd0}, waddr_nxt} : _GEN_34; // @[TensorLoad.scala 214:3:@7009.6]
  assign _GEN_37 = _T_640 ? dec_sram_offset : _GEN_35; // @[TensorLoad.scala 208:25:@6998.4]
  assign _GEN_38 = _T_640 ? dec_sram_offset : _GEN_36; // @[TensorLoad.scala 208:25:@6998.4]
  assign wmask_0_0 = tag == 3'h0; // @[TensorLoad.scala 235:26:@7037.4]
  assign wdata_0_0 = isZeroPad ? 64'h0 : io_vme_rd_data_bits; // @[TensorLoad.scala 236:25:@7039.4]
  assign wmask_0_1 = tag == 3'h1; // @[TensorLoad.scala 235:26:@7041.4]
  assign wmask_0_2 = tag == 3'h2; // @[TensorLoad.scala 235:26:@7045.4]
  assign wmask_0_3 = tag == 3'h3; // @[TensorLoad.scala 235:26:@7049.4]
  assign wmask_0_4 = tag == 3'h4; // @[TensorLoad.scala 235:26:@7053.4]
  assign wmask_0_5 = tag == 3'h5; // @[TensorLoad.scala 235:26:@7057.4]
  assign wmask_0_6 = tag == 3'h6; // @[TensorLoad.scala 235:26:@7061.4]
  assign _T_855 = {io_tensor_wr_bits_data_0_7,io_tensor_wr_bits_data_0_6,io_tensor_wr_bits_data_0_5,io_tensor_wr_bits_data_0_4,io_tensor_wr_bits_data_0_3,io_tensor_wr_bits_data_0_2,io_tensor_wr_bits_data_0_1,io_tensor_wr_bits_data_0_0}; // @[TensorLoad.scala 238:43:@7075.4]
  assign _T_863 = {io_tensor_wr_bits_data_0_15,io_tensor_wr_bits_data_0_14,io_tensor_wr_bits_data_0_13,io_tensor_wr_bits_data_0_12,io_tensor_wr_bits_data_0_11,io_tensor_wr_bits_data_0_10,io_tensor_wr_bits_data_0_9,io_tensor_wr_bits_data_0_8,_T_855}; // @[TensorLoad.scala 238:43:@7083.4]
  assign _T_915 = _T_863[63:0]; // @[TensorLoad.scala 238:58:@7087.4]
  assign _T_916 = _T_863[127:64]; // @[TensorLoad.scala 238:58:@7089.4]
  assign _T_917 = _T_863[191:128]; // @[TensorLoad.scala 238:58:@7091.4]
  assign _T_918 = _T_863[255:192]; // @[TensorLoad.scala 238:58:@7093.4]
  assign _T_919 = _T_863[319:256]; // @[TensorLoad.scala 238:58:@7095.4]
  assign _T_920 = _T_863[383:320]; // @[TensorLoad.scala 238:58:@7097.4]
  assign _T_921 = _T_863[447:384]; // @[TensorLoad.scala 238:58:@7099.4]
  assign _T_922 = _T_863[511:448]; // @[TensorLoad.scala 238:58:@7101.4]
  assign _GEN_75 = io_tensor_rd_idx_valid; // @[TensorLoad.scala 256:26:@7147.4]
  assign _T_1043 = {tensorFile_0_7_rdata_0_data,tensorFile_0_6_rdata_0_data,tensorFile_0_5_rdata_0_data,tensorFile_0_4_rdata_0_data,tensorFile_0_3_rdata_0_data,tensorFile_0_2_rdata_0_data,tensorFile_0_1_rdata_0_data,tensorFile_0_0_rdata_0_data}; // @[TensorLoad.scala 259:38:@7159.4]
  assign _T_1191 = dec_ypad_1 == 4'h0; // @[TensorLoad.scala 263:96:@7215.4]
  assign done_no_pad = _T_661 & _T_1191; // @[TensorLoad.scala 263:83:@7216.4]
  assign done_x_pad = _T_664 & _T_1191; // @[TensorLoad.scala 264:72:@7221.4]
  assign _T_1198 = _T_706 & dataCtrlDone; // @[TensorLoad.scala 265:37:@7223.4]
  assign done_y_pad = _T_1198 & yPadCtrl1_io_done; // @[TensorLoad.scala 265:52:@7224.4]
  assign _T_1199 = done_no_pad | done_x_pad; // @[TensorLoad.scala 266:26:@7225.4]
  assign io_done = _T_1199 | done_y_pad; // @[TensorLoad.scala 266:11:@7227.4]
  assign io_vme_rd_cmd_valid = state == 3'h3; // @[TensorLoad.scala 182:23:@6948.4]
  assign io_vme_rd_cmd_bits_addr = dataCtrl_io_addr; // @[TensorLoad.scala 183:27:@6949.4]
  assign io_vme_rd_cmd_bits_len = dataCtrl_io_len; // @[TensorLoad.scala 184:26:@6950.4]
  assign io_vme_rd_data_ready = state == 3'h4; // @[TensorLoad.scala 186:24:@6952.4]
  assign io_tensor_rd_data_valid = rvalid; // @[TensorLoad.scala 253:27:@7144.4]
  assign io_tensor_rd_data_bits_0_0 = _T_1043[31:0]; // @[TensorLoad.scala 259:33:@7195.4]
  assign io_tensor_rd_data_bits_0_1 = _T_1043[63:32]; // @[TensorLoad.scala 259:33:@7196.4]
  assign io_tensor_rd_data_bits_0_2 = _T_1043[95:64]; // @[TensorLoad.scala 259:33:@7197.4]
  assign io_tensor_rd_data_bits_0_3 = _T_1043[127:96]; // @[TensorLoad.scala 259:33:@7198.4]
  assign io_tensor_rd_data_bits_0_4 = _T_1043[159:128]; // @[TensorLoad.scala 259:33:@7199.4]
  assign io_tensor_rd_data_bits_0_5 = _T_1043[191:160]; // @[TensorLoad.scala 259:33:@7200.4]
  assign io_tensor_rd_data_bits_0_6 = _T_1043[223:192]; // @[TensorLoad.scala 259:33:@7201.4]
  assign io_tensor_rd_data_bits_0_7 = _T_1043[255:224]; // @[TensorLoad.scala 259:33:@7202.4]
  assign io_tensor_rd_data_bits_0_8 = _T_1043[287:256]; // @[TensorLoad.scala 259:33:@7203.4]
  assign io_tensor_rd_data_bits_0_9 = _T_1043[319:288]; // @[TensorLoad.scala 259:33:@7204.4]
  assign io_tensor_rd_data_bits_0_10 = _T_1043[351:320]; // @[TensorLoad.scala 259:33:@7205.4]
  assign io_tensor_rd_data_bits_0_11 = _T_1043[383:352]; // @[TensorLoad.scala 259:33:@7206.4]
  assign io_tensor_rd_data_bits_0_12 = _T_1043[415:384]; // @[TensorLoad.scala 259:33:@7207.4]
  assign io_tensor_rd_data_bits_0_13 = _T_1043[447:416]; // @[TensorLoad.scala 259:33:@7208.4]
  assign io_tensor_rd_data_bits_0_14 = _T_1043[479:448]; // @[TensorLoad.scala 259:33:@7209.4]
  assign io_tensor_rd_data_bits_0_15 = _T_1043[511:480]; // @[TensorLoad.scala 259:33:@7210.4]
  assign dataCtrl_clock = clock; // @[:@6743.4]
  assign dataCtrl_io_start = _T_640 & io_start; // @[TensorLoad.scala 147:21:@6878.4]
  assign dataCtrl_io_inst = io_inst; // @[TensorLoad.scala 148:20:@6879.4]
  assign dataCtrl_io_baddr = io_baddr; // @[TensorLoad.scala 149:21:@6880.4]
  assign dataCtrl_io_xinit = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[TensorLoad.scala 150:21:@6882.4]
  assign dataCtrl_io_xupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 151:23:@6884.4]
  assign dataCtrl_io_yupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 152:23:@6886.4]
  assign yPadCtrl0_clock = clock; // @[:@6747.4]
  assign yPadCtrl0_reset = reset; // @[:@6748.4]
  assign yPadCtrl0_io_start = _T_653 & io_start; // @[TensorLoad.scala 161:22:@6901.4]
  assign yPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 176:21:@6943.4]
  assign yPadCtrl1_clock = clock; // @[:@6750.4]
  assign yPadCtrl1_reset = reset; // @[:@6751.4]
  assign yPadCtrl1_io_start = _T_628 & _T_665; // @[TensorLoad.scala 163:22:@6912.4]
  assign yPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 177:21:@6944.4]
  assign xPadCtrl0_clock = clock; // @[:@6753.4]
  assign xPadCtrl0_reset = reset; // @[:@6754.4]
  assign xPadCtrl0_io_start = _T_618 & _T_686; // @[TensorLoad.scala 167:22:@6932.4]
  assign xPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 178:21:@6945.4]
  assign xPadCtrl1_clock = clock; // @[:@6756.4]
  assign xPadCtrl1_reset = reset; // @[:@6757.4]
  assign xPadCtrl1_io_start = _T_691 & _T_697; // @[TensorLoad.scala 173:22:@6942.4]
  assign xPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 179:21:@6946.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_0[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_1[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_2[initvar] = _RAND_2[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_3[initvar] = _RAND_3[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_4[initvar] = _RAND_4[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_5[initvar] = _RAND_5[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_6[initvar] = _RAND_6[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_7[initvar] = _RAND_7[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  dataCtrlDone = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  tag = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  waddr_cur = _RAND_11[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  waddr_nxt = _RAND_12[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  rvalid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  tensorFile_0_0_rdata_0_addr_pipe_0 = _RAND_14[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  tensorFile_0_1_rdata_0_addr_pipe_0 = _RAND_15[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  tensorFile_0_2_rdata_0_addr_pipe_0 = _RAND_16[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  tensorFile_0_3_rdata_0_addr_pipe_0 = _RAND_17[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  tensorFile_0_4_rdata_0_addr_pipe_0 = _RAND_18[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  tensorFile_0_5_rdata_0_addr_pipe_0 = _RAND_19[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  tensorFile_0_6_rdata_0_addr_pipe_0 = _RAND_20[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  tensorFile_0_7_rdata_0_addr_pipe_0 = _RAND_21[10:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tensorFile_0_0__T_992_en & tensorFile_0_0__T_992_mask) begin
      tensorFile_0_0[tensorFile_0_0__T_992_addr] <= tensorFile_0_0__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
    end
    if(tensorFile_0_1__T_992_en & tensorFile_0_1__T_992_mask) begin
      tensorFile_0_1[tensorFile_0_1__T_992_addr] <= tensorFile_0_1__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
    end
    if(tensorFile_0_2__T_992_en & tensorFile_0_2__T_992_mask) begin
      tensorFile_0_2[tensorFile_0_2__T_992_addr] <= tensorFile_0_2__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
    end
    if(tensorFile_0_3__T_992_en & tensorFile_0_3__T_992_mask) begin
      tensorFile_0_3[tensorFile_0_3__T_992_addr] <= tensorFile_0_3__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
    end
    if(tensorFile_0_4__T_992_en & tensorFile_0_4__T_992_mask) begin
      tensorFile_0_4[tensorFile_0_4__T_992_addr] <= tensorFile_0_4__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
    end
    if(tensorFile_0_5__T_992_en & tensorFile_0_5__T_992_mask) begin
      tensorFile_0_5[tensorFile_0_5__T_992_addr] <= tensorFile_0_5__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
    end
    if(tensorFile_0_6__T_992_en & tensorFile_0_6__T_992_mask) begin
      tensorFile_0_6[tensorFile_0_6__T_992_addr] <= tensorFile_0_6__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
    end
    if(tensorFile_0_7__T_992_en & tensorFile_0_7__T_992_mask) begin
      tensorFile_0_7[tensorFile_0_7__T_992_addr] <= tensorFile_0_7__T_992_data; // @[TensorLoad.scala 222:16:@7025.4]
    end
    if (reset) begin
      dataCtrlDone <= 1'h0;
    end else begin
      if (_T_640) begin
        dataCtrlDone <= 1'h0;
      end else begin
        if (_T_648) begin
          dataCtrlDone <= 1'h1;
        end
      end
    end
    if (_T_712) begin
      tag <= 3'h0;
    end else begin
      if (_T_715) begin
        tag <= _T_718;
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_614) begin
        if (io_start) begin
          if (_T_616) begin
            state <= 3'h1;
          end else begin
            if (_T_618) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end
      end else begin
        if (_T_619) begin
          if (yPadCtrl0_io_done) begin
            if (_T_618) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end else begin
          if (_T_622) begin
            if (xPadCtrl0_io_done) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_623) begin
              if (io_vme_rd_cmd_ready) begin
                state <= 3'h4;
              end
            end else begin
              if (_T_624) begin
                if (io_vme_rd_data_valid) begin
                  if (dataCtrl_io_done) begin
                    if (_T_626) begin
                      state <= 3'h5;
                    end else begin
                      if (_T_628) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end
                  end else begin
                    if (dataCtrl_io_stride) begin
                      if (_T_626) begin
                        state <= 3'h5;
                      end else begin
                        if (_T_618) begin
                          state <= 3'h2;
                        end else begin
                          state <= 3'h3;
                        end
                      end
                    end else begin
                      if (dataCtrl_io_split) begin
                        state <= 3'h3;
                      end
                    end
                  end
                end
              end else begin
                if (_T_633) begin
                  if (xPadCtrl1_io_done) begin
                    if (dataCtrlDone) begin
                      if (_T_628) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end else begin
                      if (_T_618) begin
                        state <= 3'h2;
                      end else begin
                        state <= 3'h3;
                      end
                    end
                  end
                end else begin
                  if (_T_638) begin
                    if (_T_639) begin
                      state <= 3'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    waddr_cur <= _GEN_37[10:0];
    waddr_nxt <= _GEN_38[10:0];
    rvalid <= io_tensor_rd_idx_valid;
    if (_GEN_75) begin
      tensorFile_0_0_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_1_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_2_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_3_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_4_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_5_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_6_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_7_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
  end
endmodule
module MAC( // @[:@7229.2]
  input         clock, // @[:@7230.4]
  input  [7:0]  io_a, // @[:@7232.4]
  input  [7:0]  io_b, // @[:@7232.4]
  input         io_c, // @[:@7232.4]
  output [16:0] io_y // @[:@7232.4]
);
  reg [7:0] rA; // @[TensorGemm.scala 39:19:@7236.4]
  reg [31:0] _RAND_0;
  reg [7:0] rB; // @[TensorGemm.scala 40:19:@7238.4]
  reg [31:0] _RAND_1;
  reg  rC; // @[TensorGemm.scala 41:19:@7240.4]
  reg [31:0] _RAND_2;
  wire [15:0] mult; // @[TensorGemm.scala 43:14:@7242.4]
  wire [15:0] _GEN_0; // @[TensorGemm.scala 44:13:@7244.4]
  assign mult = $signed(rA) * $signed(rB); // @[TensorGemm.scala 43:14:@7242.4]
  assign _GEN_0 = {16{rC}}; // @[TensorGemm.scala 44:13:@7244.4]
  assign io_y = $signed(_GEN_0) + $signed(mult); // @[TensorGemm.scala 46:8:@7246.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rA = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rB = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rC = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    rA <= io_a;
    rB <= io_b;
    rC <= io_c;
  end
endmodule
module PipeAdder( // @[:@7533.2]
  input         clock, // @[:@7534.4]
  input  [16:0] io_a, // @[:@7536.4]
  input  [16:0] io_b, // @[:@7536.4]
  output [17:0] io_y // @[:@7536.4]
);
  reg [16:0] rA; // @[TensorGemm.scala 61:19:@7539.4]
  reg [31:0] _RAND_0;
  reg [16:0] rB; // @[TensorGemm.scala 62:19:@7541.4]
  reg [31:0] _RAND_1;
  assign io_y = $signed(rA) + $signed(rB); // @[TensorGemm.scala 64:8:@7545.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rA = _RAND_0[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rB = _RAND_1[16:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    rA <= io_a;
    rB <= io_b;
  end
endmodule
module Adder( // @[:@7645.2]
  input  [17:0] io_a, // @[:@7648.4]
  input  [17:0] io_b, // @[:@7648.4]
  output [18:0] io_y // @[:@7648.4]
);
  assign io_y = $signed(io_a) + $signed(io_b); // @[TensorGemm.scala 85:8:@7657.4]
endmodule
module Adder_4( // @[:@7701.2]
  input  [18:0] io_a, // @[:@7704.4]
  input  [18:0] io_b, // @[:@7704.4]
  output [19:0] io_y // @[:@7704.4]
);
  assign io_y = $signed(io_a) + $signed(io_b); // @[TensorGemm.scala 85:8:@7713.4]
endmodule
module Adder_6( // @[:@7729.2]
  input  [19:0] io_a, // @[:@7732.4]
  input  [19:0] io_b, // @[:@7732.4]
  output [20:0] io_y // @[:@7732.4]
);
  assign io_y = $signed(io_a) + $signed(io_b); // @[TensorGemm.scala 85:8:@7741.4]
endmodule
module DotProduct( // @[:@7743.2]
  input         clock, // @[:@7744.4]
  input  [7:0]  io_a_0, // @[:@7746.4]
  input  [7:0]  io_a_1, // @[:@7746.4]
  input  [7:0]  io_a_2, // @[:@7746.4]
  input  [7:0]  io_a_3, // @[:@7746.4]
  input  [7:0]  io_a_4, // @[:@7746.4]
  input  [7:0]  io_a_5, // @[:@7746.4]
  input  [7:0]  io_a_6, // @[:@7746.4]
  input  [7:0]  io_a_7, // @[:@7746.4]
  input  [7:0]  io_a_8, // @[:@7746.4]
  input  [7:0]  io_a_9, // @[:@7746.4]
  input  [7:0]  io_a_10, // @[:@7746.4]
  input  [7:0]  io_a_11, // @[:@7746.4]
  input  [7:0]  io_a_12, // @[:@7746.4]
  input  [7:0]  io_a_13, // @[:@7746.4]
  input  [7:0]  io_a_14, // @[:@7746.4]
  input  [7:0]  io_a_15, // @[:@7746.4]
  input  [7:0]  io_b_0, // @[:@7746.4]
  input  [7:0]  io_b_1, // @[:@7746.4]
  input  [7:0]  io_b_2, // @[:@7746.4]
  input  [7:0]  io_b_3, // @[:@7746.4]
  input  [7:0]  io_b_4, // @[:@7746.4]
  input  [7:0]  io_b_5, // @[:@7746.4]
  input  [7:0]  io_b_6, // @[:@7746.4]
  input  [7:0]  io_b_7, // @[:@7746.4]
  input  [7:0]  io_b_8, // @[:@7746.4]
  input  [7:0]  io_b_9, // @[:@7746.4]
  input  [7:0]  io_b_10, // @[:@7746.4]
  input  [7:0]  io_b_11, // @[:@7746.4]
  input  [7:0]  io_b_12, // @[:@7746.4]
  input  [7:0]  io_b_13, // @[:@7746.4]
  input  [7:0]  io_b_14, // @[:@7746.4]
  input  [7:0]  io_b_15, // @[:@7746.4]
  output [20:0] io_y // @[:@7746.4]
);
  wire  m_0_clock; // @[TensorGemm.scala 103:32:@7748.4]
  wire [7:0] m_0_io_a; // @[TensorGemm.scala 103:32:@7748.4]
  wire [7:0] m_0_io_b; // @[TensorGemm.scala 103:32:@7748.4]
  wire  m_0_io_c; // @[TensorGemm.scala 103:32:@7748.4]
  wire [16:0] m_0_io_y; // @[TensorGemm.scala 103:32:@7748.4]
  wire  m_1_clock; // @[TensorGemm.scala 103:32:@7751.4]
  wire [7:0] m_1_io_a; // @[TensorGemm.scala 103:32:@7751.4]
  wire [7:0] m_1_io_b; // @[TensorGemm.scala 103:32:@7751.4]
  wire  m_1_io_c; // @[TensorGemm.scala 103:32:@7751.4]
  wire [16:0] m_1_io_y; // @[TensorGemm.scala 103:32:@7751.4]
  wire  m_2_clock; // @[TensorGemm.scala 103:32:@7754.4]
  wire [7:0] m_2_io_a; // @[TensorGemm.scala 103:32:@7754.4]
  wire [7:0] m_2_io_b; // @[TensorGemm.scala 103:32:@7754.4]
  wire  m_2_io_c; // @[TensorGemm.scala 103:32:@7754.4]
  wire [16:0] m_2_io_y; // @[TensorGemm.scala 103:32:@7754.4]
  wire  m_3_clock; // @[TensorGemm.scala 103:32:@7757.4]
  wire [7:0] m_3_io_a; // @[TensorGemm.scala 103:32:@7757.4]
  wire [7:0] m_3_io_b; // @[TensorGemm.scala 103:32:@7757.4]
  wire  m_3_io_c; // @[TensorGemm.scala 103:32:@7757.4]
  wire [16:0] m_3_io_y; // @[TensorGemm.scala 103:32:@7757.4]
  wire  m_4_clock; // @[TensorGemm.scala 103:32:@7760.4]
  wire [7:0] m_4_io_a; // @[TensorGemm.scala 103:32:@7760.4]
  wire [7:0] m_4_io_b; // @[TensorGemm.scala 103:32:@7760.4]
  wire  m_4_io_c; // @[TensorGemm.scala 103:32:@7760.4]
  wire [16:0] m_4_io_y; // @[TensorGemm.scala 103:32:@7760.4]
  wire  m_5_clock; // @[TensorGemm.scala 103:32:@7763.4]
  wire [7:0] m_5_io_a; // @[TensorGemm.scala 103:32:@7763.4]
  wire [7:0] m_5_io_b; // @[TensorGemm.scala 103:32:@7763.4]
  wire  m_5_io_c; // @[TensorGemm.scala 103:32:@7763.4]
  wire [16:0] m_5_io_y; // @[TensorGemm.scala 103:32:@7763.4]
  wire  m_6_clock; // @[TensorGemm.scala 103:32:@7766.4]
  wire [7:0] m_6_io_a; // @[TensorGemm.scala 103:32:@7766.4]
  wire [7:0] m_6_io_b; // @[TensorGemm.scala 103:32:@7766.4]
  wire  m_6_io_c; // @[TensorGemm.scala 103:32:@7766.4]
  wire [16:0] m_6_io_y; // @[TensorGemm.scala 103:32:@7766.4]
  wire  m_7_clock; // @[TensorGemm.scala 103:32:@7769.4]
  wire [7:0] m_7_io_a; // @[TensorGemm.scala 103:32:@7769.4]
  wire [7:0] m_7_io_b; // @[TensorGemm.scala 103:32:@7769.4]
  wire  m_7_io_c; // @[TensorGemm.scala 103:32:@7769.4]
  wire [16:0] m_7_io_y; // @[TensorGemm.scala 103:32:@7769.4]
  wire  m_8_clock; // @[TensorGemm.scala 103:32:@7772.4]
  wire [7:0] m_8_io_a; // @[TensorGemm.scala 103:32:@7772.4]
  wire [7:0] m_8_io_b; // @[TensorGemm.scala 103:32:@7772.4]
  wire  m_8_io_c; // @[TensorGemm.scala 103:32:@7772.4]
  wire [16:0] m_8_io_y; // @[TensorGemm.scala 103:32:@7772.4]
  wire  m_9_clock; // @[TensorGemm.scala 103:32:@7775.4]
  wire [7:0] m_9_io_a; // @[TensorGemm.scala 103:32:@7775.4]
  wire [7:0] m_9_io_b; // @[TensorGemm.scala 103:32:@7775.4]
  wire  m_9_io_c; // @[TensorGemm.scala 103:32:@7775.4]
  wire [16:0] m_9_io_y; // @[TensorGemm.scala 103:32:@7775.4]
  wire  m_10_clock; // @[TensorGemm.scala 103:32:@7778.4]
  wire [7:0] m_10_io_a; // @[TensorGemm.scala 103:32:@7778.4]
  wire [7:0] m_10_io_b; // @[TensorGemm.scala 103:32:@7778.4]
  wire  m_10_io_c; // @[TensorGemm.scala 103:32:@7778.4]
  wire [16:0] m_10_io_y; // @[TensorGemm.scala 103:32:@7778.4]
  wire  m_11_clock; // @[TensorGemm.scala 103:32:@7781.4]
  wire [7:0] m_11_io_a; // @[TensorGemm.scala 103:32:@7781.4]
  wire [7:0] m_11_io_b; // @[TensorGemm.scala 103:32:@7781.4]
  wire  m_11_io_c; // @[TensorGemm.scala 103:32:@7781.4]
  wire [16:0] m_11_io_y; // @[TensorGemm.scala 103:32:@7781.4]
  wire  m_12_clock; // @[TensorGemm.scala 103:32:@7784.4]
  wire [7:0] m_12_io_a; // @[TensorGemm.scala 103:32:@7784.4]
  wire [7:0] m_12_io_b; // @[TensorGemm.scala 103:32:@7784.4]
  wire  m_12_io_c; // @[TensorGemm.scala 103:32:@7784.4]
  wire [16:0] m_12_io_y; // @[TensorGemm.scala 103:32:@7784.4]
  wire  m_13_clock; // @[TensorGemm.scala 103:32:@7787.4]
  wire [7:0] m_13_io_a; // @[TensorGemm.scala 103:32:@7787.4]
  wire [7:0] m_13_io_b; // @[TensorGemm.scala 103:32:@7787.4]
  wire  m_13_io_c; // @[TensorGemm.scala 103:32:@7787.4]
  wire [16:0] m_13_io_y; // @[TensorGemm.scala 103:32:@7787.4]
  wire  m_14_clock; // @[TensorGemm.scala 103:32:@7790.4]
  wire [7:0] m_14_io_a; // @[TensorGemm.scala 103:32:@7790.4]
  wire [7:0] m_14_io_b; // @[TensorGemm.scala 103:32:@7790.4]
  wire  m_14_io_c; // @[TensorGemm.scala 103:32:@7790.4]
  wire [16:0] m_14_io_y; // @[TensorGemm.scala 103:32:@7790.4]
  wire  m_15_clock; // @[TensorGemm.scala 103:32:@7793.4]
  wire [7:0] m_15_io_a; // @[TensorGemm.scala 103:32:@7793.4]
  wire [7:0] m_15_io_b; // @[TensorGemm.scala 103:32:@7793.4]
  wire  m_15_io_c; // @[TensorGemm.scala 103:32:@7793.4]
  wire [16:0] m_15_io_y; // @[TensorGemm.scala 103:32:@7793.4]
  wire  a_0_0_clock; // @[TensorGemm.scala 108:17:@7796.4]
  wire [16:0] a_0_0_io_a; // @[TensorGemm.scala 108:17:@7796.4]
  wire [16:0] a_0_0_io_b; // @[TensorGemm.scala 108:17:@7796.4]
  wire [17:0] a_0_0_io_y; // @[TensorGemm.scala 108:17:@7796.4]
  wire  a_0_1_clock; // @[TensorGemm.scala 108:17:@7799.4]
  wire [16:0] a_0_1_io_a; // @[TensorGemm.scala 108:17:@7799.4]
  wire [16:0] a_0_1_io_b; // @[TensorGemm.scala 108:17:@7799.4]
  wire [17:0] a_0_1_io_y; // @[TensorGemm.scala 108:17:@7799.4]
  wire  a_0_2_clock; // @[TensorGemm.scala 108:17:@7802.4]
  wire [16:0] a_0_2_io_a; // @[TensorGemm.scala 108:17:@7802.4]
  wire [16:0] a_0_2_io_b; // @[TensorGemm.scala 108:17:@7802.4]
  wire [17:0] a_0_2_io_y; // @[TensorGemm.scala 108:17:@7802.4]
  wire  a_0_3_clock; // @[TensorGemm.scala 108:17:@7805.4]
  wire [16:0] a_0_3_io_a; // @[TensorGemm.scala 108:17:@7805.4]
  wire [16:0] a_0_3_io_b; // @[TensorGemm.scala 108:17:@7805.4]
  wire [17:0] a_0_3_io_y; // @[TensorGemm.scala 108:17:@7805.4]
  wire  a_0_4_clock; // @[TensorGemm.scala 108:17:@7808.4]
  wire [16:0] a_0_4_io_a; // @[TensorGemm.scala 108:17:@7808.4]
  wire [16:0] a_0_4_io_b; // @[TensorGemm.scala 108:17:@7808.4]
  wire [17:0] a_0_4_io_y; // @[TensorGemm.scala 108:17:@7808.4]
  wire  a_0_5_clock; // @[TensorGemm.scala 108:17:@7811.4]
  wire [16:0] a_0_5_io_a; // @[TensorGemm.scala 108:17:@7811.4]
  wire [16:0] a_0_5_io_b; // @[TensorGemm.scala 108:17:@7811.4]
  wire [17:0] a_0_5_io_y; // @[TensorGemm.scala 108:17:@7811.4]
  wire  a_0_6_clock; // @[TensorGemm.scala 108:17:@7814.4]
  wire [16:0] a_0_6_io_a; // @[TensorGemm.scala 108:17:@7814.4]
  wire [16:0] a_0_6_io_b; // @[TensorGemm.scala 108:17:@7814.4]
  wire [17:0] a_0_6_io_y; // @[TensorGemm.scala 108:17:@7814.4]
  wire  a_0_7_clock; // @[TensorGemm.scala 108:17:@7817.4]
  wire [16:0] a_0_7_io_a; // @[TensorGemm.scala 108:17:@7817.4]
  wire [16:0] a_0_7_io_b; // @[TensorGemm.scala 108:17:@7817.4]
  wire [17:0] a_0_7_io_y; // @[TensorGemm.scala 108:17:@7817.4]
  wire [17:0] a_1_0_io_a; // @[TensorGemm.scala 110:17:@7820.4]
  wire [17:0] a_1_0_io_b; // @[TensorGemm.scala 110:17:@7820.4]
  wire [18:0] a_1_0_io_y; // @[TensorGemm.scala 110:17:@7820.4]
  wire [17:0] a_1_1_io_a; // @[TensorGemm.scala 110:17:@7823.4]
  wire [17:0] a_1_1_io_b; // @[TensorGemm.scala 110:17:@7823.4]
  wire [18:0] a_1_1_io_y; // @[TensorGemm.scala 110:17:@7823.4]
  wire [17:0] a_1_2_io_a; // @[TensorGemm.scala 110:17:@7826.4]
  wire [17:0] a_1_2_io_b; // @[TensorGemm.scala 110:17:@7826.4]
  wire [18:0] a_1_2_io_y; // @[TensorGemm.scala 110:17:@7826.4]
  wire [17:0] a_1_3_io_a; // @[TensorGemm.scala 110:17:@7829.4]
  wire [17:0] a_1_3_io_b; // @[TensorGemm.scala 110:17:@7829.4]
  wire [18:0] a_1_3_io_y; // @[TensorGemm.scala 110:17:@7829.4]
  wire [18:0] a_2_0_io_a; // @[TensorGemm.scala 110:17:@7832.4]
  wire [18:0] a_2_0_io_b; // @[TensorGemm.scala 110:17:@7832.4]
  wire [19:0] a_2_0_io_y; // @[TensorGemm.scala 110:17:@7832.4]
  wire [18:0] a_2_1_io_a; // @[TensorGemm.scala 110:17:@7835.4]
  wire [18:0] a_2_1_io_b; // @[TensorGemm.scala 110:17:@7835.4]
  wire [19:0] a_2_1_io_y; // @[TensorGemm.scala 110:17:@7835.4]
  wire [19:0] a_3_0_io_a; // @[TensorGemm.scala 110:17:@7838.4]
  wire [19:0] a_3_0_io_b; // @[TensorGemm.scala 110:17:@7838.4]
  wire [20:0] a_3_0_io_y; // @[TensorGemm.scala 110:17:@7838.4]
  MAC m_0 ( // @[TensorGemm.scala 103:32:@7748.4]
    .clock(m_0_clock),
    .io_a(m_0_io_a),
    .io_b(m_0_io_b),
    .io_c(m_0_io_c),
    .io_y(m_0_io_y)
  );
  MAC m_1 ( // @[TensorGemm.scala 103:32:@7751.4]
    .clock(m_1_clock),
    .io_a(m_1_io_a),
    .io_b(m_1_io_b),
    .io_c(m_1_io_c),
    .io_y(m_1_io_y)
  );
  MAC m_2 ( // @[TensorGemm.scala 103:32:@7754.4]
    .clock(m_2_clock),
    .io_a(m_2_io_a),
    .io_b(m_2_io_b),
    .io_c(m_2_io_c),
    .io_y(m_2_io_y)
  );
  MAC m_3 ( // @[TensorGemm.scala 103:32:@7757.4]
    .clock(m_3_clock),
    .io_a(m_3_io_a),
    .io_b(m_3_io_b),
    .io_c(m_3_io_c),
    .io_y(m_3_io_y)
  );
  MAC m_4 ( // @[TensorGemm.scala 103:32:@7760.4]
    .clock(m_4_clock),
    .io_a(m_4_io_a),
    .io_b(m_4_io_b),
    .io_c(m_4_io_c),
    .io_y(m_4_io_y)
  );
  MAC m_5 ( // @[TensorGemm.scala 103:32:@7763.4]
    .clock(m_5_clock),
    .io_a(m_5_io_a),
    .io_b(m_5_io_b),
    .io_c(m_5_io_c),
    .io_y(m_5_io_y)
  );
  MAC m_6 ( // @[TensorGemm.scala 103:32:@7766.4]
    .clock(m_6_clock),
    .io_a(m_6_io_a),
    .io_b(m_6_io_b),
    .io_c(m_6_io_c),
    .io_y(m_6_io_y)
  );
  MAC m_7 ( // @[TensorGemm.scala 103:32:@7769.4]
    .clock(m_7_clock),
    .io_a(m_7_io_a),
    .io_b(m_7_io_b),
    .io_c(m_7_io_c),
    .io_y(m_7_io_y)
  );
  MAC m_8 ( // @[TensorGemm.scala 103:32:@7772.4]
    .clock(m_8_clock),
    .io_a(m_8_io_a),
    .io_b(m_8_io_b),
    .io_c(m_8_io_c),
    .io_y(m_8_io_y)
  );
  MAC m_9 ( // @[TensorGemm.scala 103:32:@7775.4]
    .clock(m_9_clock),
    .io_a(m_9_io_a),
    .io_b(m_9_io_b),
    .io_c(m_9_io_c),
    .io_y(m_9_io_y)
  );
  MAC m_10 ( // @[TensorGemm.scala 103:32:@7778.4]
    .clock(m_10_clock),
    .io_a(m_10_io_a),
    .io_b(m_10_io_b),
    .io_c(m_10_io_c),
    .io_y(m_10_io_y)
  );
  MAC m_11 ( // @[TensorGemm.scala 103:32:@7781.4]
    .clock(m_11_clock),
    .io_a(m_11_io_a),
    .io_b(m_11_io_b),
    .io_c(m_11_io_c),
    .io_y(m_11_io_y)
  );
  MAC m_12 ( // @[TensorGemm.scala 103:32:@7784.4]
    .clock(m_12_clock),
    .io_a(m_12_io_a),
    .io_b(m_12_io_b),
    .io_c(m_12_io_c),
    .io_y(m_12_io_y)
  );
  MAC m_13 ( // @[TensorGemm.scala 103:32:@7787.4]
    .clock(m_13_clock),
    .io_a(m_13_io_a),
    .io_b(m_13_io_b),
    .io_c(m_13_io_c),
    .io_y(m_13_io_y)
  );
  MAC m_14 ( // @[TensorGemm.scala 103:32:@7790.4]
    .clock(m_14_clock),
    .io_a(m_14_io_a),
    .io_b(m_14_io_b),
    .io_c(m_14_io_c),
    .io_y(m_14_io_y)
  );
  MAC m_15 ( // @[TensorGemm.scala 103:32:@7793.4]
    .clock(m_15_clock),
    .io_a(m_15_io_a),
    .io_b(m_15_io_b),
    .io_c(m_15_io_c),
    .io_y(m_15_io_y)
  );
  PipeAdder a_0_0 ( // @[TensorGemm.scala 108:17:@7796.4]
    .clock(a_0_0_clock),
    .io_a(a_0_0_io_a),
    .io_b(a_0_0_io_b),
    .io_y(a_0_0_io_y)
  );
  PipeAdder a_0_1 ( // @[TensorGemm.scala 108:17:@7799.4]
    .clock(a_0_1_clock),
    .io_a(a_0_1_io_a),
    .io_b(a_0_1_io_b),
    .io_y(a_0_1_io_y)
  );
  PipeAdder a_0_2 ( // @[TensorGemm.scala 108:17:@7802.4]
    .clock(a_0_2_clock),
    .io_a(a_0_2_io_a),
    .io_b(a_0_2_io_b),
    .io_y(a_0_2_io_y)
  );
  PipeAdder a_0_3 ( // @[TensorGemm.scala 108:17:@7805.4]
    .clock(a_0_3_clock),
    .io_a(a_0_3_io_a),
    .io_b(a_0_3_io_b),
    .io_y(a_0_3_io_y)
  );
  PipeAdder a_0_4 ( // @[TensorGemm.scala 108:17:@7808.4]
    .clock(a_0_4_clock),
    .io_a(a_0_4_io_a),
    .io_b(a_0_4_io_b),
    .io_y(a_0_4_io_y)
  );
  PipeAdder a_0_5 ( // @[TensorGemm.scala 108:17:@7811.4]
    .clock(a_0_5_clock),
    .io_a(a_0_5_io_a),
    .io_b(a_0_5_io_b),
    .io_y(a_0_5_io_y)
  );
  PipeAdder a_0_6 ( // @[TensorGemm.scala 108:17:@7814.4]
    .clock(a_0_6_clock),
    .io_a(a_0_6_io_a),
    .io_b(a_0_6_io_b),
    .io_y(a_0_6_io_y)
  );
  PipeAdder a_0_7 ( // @[TensorGemm.scala 108:17:@7817.4]
    .clock(a_0_7_clock),
    .io_a(a_0_7_io_a),
    .io_b(a_0_7_io_b),
    .io_y(a_0_7_io_y)
  );
  Adder a_1_0 ( // @[TensorGemm.scala 110:17:@7820.4]
    .io_a(a_1_0_io_a),
    .io_b(a_1_0_io_b),
    .io_y(a_1_0_io_y)
  );
  Adder a_1_1 ( // @[TensorGemm.scala 110:17:@7823.4]
    .io_a(a_1_1_io_a),
    .io_b(a_1_1_io_b),
    .io_y(a_1_1_io_y)
  );
  Adder a_1_2 ( // @[TensorGemm.scala 110:17:@7826.4]
    .io_a(a_1_2_io_a),
    .io_b(a_1_2_io_b),
    .io_y(a_1_2_io_y)
  );
  Adder a_1_3 ( // @[TensorGemm.scala 110:17:@7829.4]
    .io_a(a_1_3_io_a),
    .io_b(a_1_3_io_b),
    .io_y(a_1_3_io_y)
  );
  Adder_4 a_2_0 ( // @[TensorGemm.scala 110:17:@7832.4]
    .io_a(a_2_0_io_a),
    .io_b(a_2_0_io_b),
    .io_y(a_2_0_io_y)
  );
  Adder_4 a_2_1 ( // @[TensorGemm.scala 110:17:@7835.4]
    .io_a(a_2_1_io_a),
    .io_b(a_2_1_io_b),
    .io_y(a_2_1_io_y)
  );
  Adder_6 a_3_0 ( // @[TensorGemm.scala 110:17:@7838.4]
    .io_a(a_3_0_io_a),
    .io_b(a_3_0_io_b),
    .io_y(a_3_0_io_y)
  );
  assign io_y = a_3_0_io_y; // @[TensorGemm.scala 134:8:@7919.4]
  assign m_0_clock = clock; // @[:@7749.4]
  assign m_0_io_a = io_a_0; // @[TensorGemm.scala 114:15:@7841.4]
  assign m_0_io_b = io_b_0; // @[TensorGemm.scala 115:15:@7842.4]
  assign m_0_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7843.4]
  assign m_1_clock = clock; // @[:@7752.4]
  assign m_1_io_a = io_a_1; // @[TensorGemm.scala 114:15:@7844.4]
  assign m_1_io_b = io_b_1; // @[TensorGemm.scala 115:15:@7845.4]
  assign m_1_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7846.4]
  assign m_2_clock = clock; // @[:@7755.4]
  assign m_2_io_a = io_a_2; // @[TensorGemm.scala 114:15:@7847.4]
  assign m_2_io_b = io_b_2; // @[TensorGemm.scala 115:15:@7848.4]
  assign m_2_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7849.4]
  assign m_3_clock = clock; // @[:@7758.4]
  assign m_3_io_a = io_a_3; // @[TensorGemm.scala 114:15:@7850.4]
  assign m_3_io_b = io_b_3; // @[TensorGemm.scala 115:15:@7851.4]
  assign m_3_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7852.4]
  assign m_4_clock = clock; // @[:@7761.4]
  assign m_4_io_a = io_a_4; // @[TensorGemm.scala 114:15:@7853.4]
  assign m_4_io_b = io_b_4; // @[TensorGemm.scala 115:15:@7854.4]
  assign m_4_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7855.4]
  assign m_5_clock = clock; // @[:@7764.4]
  assign m_5_io_a = io_a_5; // @[TensorGemm.scala 114:15:@7856.4]
  assign m_5_io_b = io_b_5; // @[TensorGemm.scala 115:15:@7857.4]
  assign m_5_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7858.4]
  assign m_6_clock = clock; // @[:@7767.4]
  assign m_6_io_a = io_a_6; // @[TensorGemm.scala 114:15:@7859.4]
  assign m_6_io_b = io_b_6; // @[TensorGemm.scala 115:15:@7860.4]
  assign m_6_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7861.4]
  assign m_7_clock = clock; // @[:@7770.4]
  assign m_7_io_a = io_a_7; // @[TensorGemm.scala 114:15:@7862.4]
  assign m_7_io_b = io_b_7; // @[TensorGemm.scala 115:15:@7863.4]
  assign m_7_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7864.4]
  assign m_8_clock = clock; // @[:@7773.4]
  assign m_8_io_a = io_a_8; // @[TensorGemm.scala 114:15:@7865.4]
  assign m_8_io_b = io_b_8; // @[TensorGemm.scala 115:15:@7866.4]
  assign m_8_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7867.4]
  assign m_9_clock = clock; // @[:@7776.4]
  assign m_9_io_a = io_a_9; // @[TensorGemm.scala 114:15:@7868.4]
  assign m_9_io_b = io_b_9; // @[TensorGemm.scala 115:15:@7869.4]
  assign m_9_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7870.4]
  assign m_10_clock = clock; // @[:@7779.4]
  assign m_10_io_a = io_a_10; // @[TensorGemm.scala 114:15:@7871.4]
  assign m_10_io_b = io_b_10; // @[TensorGemm.scala 115:15:@7872.4]
  assign m_10_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7873.4]
  assign m_11_clock = clock; // @[:@7782.4]
  assign m_11_io_a = io_a_11; // @[TensorGemm.scala 114:15:@7874.4]
  assign m_11_io_b = io_b_11; // @[TensorGemm.scala 115:15:@7875.4]
  assign m_11_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7876.4]
  assign m_12_clock = clock; // @[:@7785.4]
  assign m_12_io_a = io_a_12; // @[TensorGemm.scala 114:15:@7877.4]
  assign m_12_io_b = io_b_12; // @[TensorGemm.scala 115:15:@7878.4]
  assign m_12_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7879.4]
  assign m_13_clock = clock; // @[:@7788.4]
  assign m_13_io_a = io_a_13; // @[TensorGemm.scala 114:15:@7880.4]
  assign m_13_io_b = io_b_13; // @[TensorGemm.scala 115:15:@7881.4]
  assign m_13_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7882.4]
  assign m_14_clock = clock; // @[:@7791.4]
  assign m_14_io_a = io_a_14; // @[TensorGemm.scala 114:15:@7883.4]
  assign m_14_io_b = io_b_14; // @[TensorGemm.scala 115:15:@7884.4]
  assign m_14_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7885.4]
  assign m_15_clock = clock; // @[:@7794.4]
  assign m_15_io_a = io_a_15; // @[TensorGemm.scala 114:15:@7886.4]
  assign m_15_io_b = io_b_15; // @[TensorGemm.scala 115:15:@7887.4]
  assign m_15_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@7888.4]
  assign a_0_0_clock = clock; // @[:@7797.4]
  assign a_0_0_io_a = m_0_io_y; // @[TensorGemm.scala 124:22:@7889.4]
  assign a_0_0_io_b = m_1_io_y; // @[TensorGemm.scala 125:22:@7890.4]
  assign a_0_1_clock = clock; // @[:@7800.4]
  assign a_0_1_io_a = m_2_io_y; // @[TensorGemm.scala 124:22:@7891.4]
  assign a_0_1_io_b = m_3_io_y; // @[TensorGemm.scala 125:22:@7892.4]
  assign a_0_2_clock = clock; // @[:@7803.4]
  assign a_0_2_io_a = m_4_io_y; // @[TensorGemm.scala 124:22:@7893.4]
  assign a_0_2_io_b = m_5_io_y; // @[TensorGemm.scala 125:22:@7894.4]
  assign a_0_3_clock = clock; // @[:@7806.4]
  assign a_0_3_io_a = m_6_io_y; // @[TensorGemm.scala 124:22:@7895.4]
  assign a_0_3_io_b = m_7_io_y; // @[TensorGemm.scala 125:22:@7896.4]
  assign a_0_4_clock = clock; // @[:@7809.4]
  assign a_0_4_io_a = m_8_io_y; // @[TensorGemm.scala 124:22:@7897.4]
  assign a_0_4_io_b = m_9_io_y; // @[TensorGemm.scala 125:22:@7898.4]
  assign a_0_5_clock = clock; // @[:@7812.4]
  assign a_0_5_io_a = m_10_io_y; // @[TensorGemm.scala 124:22:@7899.4]
  assign a_0_5_io_b = m_11_io_y; // @[TensorGemm.scala 125:22:@7900.4]
  assign a_0_6_clock = clock; // @[:@7815.4]
  assign a_0_6_io_a = m_12_io_y; // @[TensorGemm.scala 124:22:@7901.4]
  assign a_0_6_io_b = m_13_io_y; // @[TensorGemm.scala 125:22:@7902.4]
  assign a_0_7_clock = clock; // @[:@7818.4]
  assign a_0_7_io_a = m_14_io_y; // @[TensorGemm.scala 124:22:@7903.4]
  assign a_0_7_io_b = m_15_io_y; // @[TensorGemm.scala 125:22:@7904.4]
  assign a_1_0_io_a = a_0_0_io_y; // @[TensorGemm.scala 127:22:@7905.4]
  assign a_1_0_io_b = a_0_1_io_y; // @[TensorGemm.scala 128:22:@7906.4]
  assign a_1_1_io_a = a_0_2_io_y; // @[TensorGemm.scala 127:22:@7907.4]
  assign a_1_1_io_b = a_0_3_io_y; // @[TensorGemm.scala 128:22:@7908.4]
  assign a_1_2_io_a = a_0_4_io_y; // @[TensorGemm.scala 127:22:@7909.4]
  assign a_1_2_io_b = a_0_5_io_y; // @[TensorGemm.scala 128:22:@7910.4]
  assign a_1_3_io_a = a_0_6_io_y; // @[TensorGemm.scala 127:22:@7911.4]
  assign a_1_3_io_b = a_0_7_io_y; // @[TensorGemm.scala 128:22:@7912.4]
  assign a_2_0_io_a = a_1_0_io_y; // @[TensorGemm.scala 127:22:@7913.4]
  assign a_2_0_io_b = a_1_1_io_y; // @[TensorGemm.scala 128:22:@7914.4]
  assign a_2_1_io_a = a_1_2_io_y; // @[TensorGemm.scala 127:22:@7915.4]
  assign a_2_1_io_b = a_1_3_io_y; // @[TensorGemm.scala 128:22:@7916.4]
  assign a_3_0_io_a = a_2_0_io_y; // @[TensorGemm.scala 127:22:@7917.4]
  assign a_3_0_io_b = a_2_1_io_y; // @[TensorGemm.scala 128:22:@7918.4]
endmodule
module Pipe( // @[:@18301.2]
  input         clock, // @[:@18302.4]
  input         reset, // @[:@18303.4]
  input         io_enq_valid, // @[:@18304.4]
  input  [31:0] io_enq_bits, // @[:@18304.4]
  output        io_deq_valid, // @[:@18304.4]
  output [31:0] io_deq_bits // @[:@18304.4]
);
  reg  _T_19; // @[Valid.scala 48:22:@18306.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_21; // @[Reg.scala 11:16:@18308.4]
  reg [31:0] _RAND_1;
  reg  _T_24; // @[Valid.scala 48:22:@18312.4]
  reg [31:0] _RAND_2;
  reg [31:0] _T_26; // @[Reg.scala 11:16:@18314.4]
  reg [31:0] _RAND_3;
  assign io_deq_valid = _T_24; // @[Valid.scala 70:10:@18322.4]
  assign io_deq_bits = _T_26; // @[Valid.scala 70:10:@18321.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_21 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_24 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_26 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      _T_19 <= io_enq_valid;
    end
    if (io_enq_valid) begin
      _T_21 <= io_enq_bits;
    end
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_19;
    end
    if (_T_19) begin
      _T_26 <= _T_21;
    end
  end
endmodule
module MatrixVectorMultiplication( // @[:@18669.2]
  input         clock, // @[:@18670.4]
  input         reset, // @[:@18671.4]
  input         io_reset, // @[:@18672.4]
  input         io_inp_data_valid, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_0, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_1, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_2, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_3, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_4, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_5, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_6, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_7, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_8, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_9, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_10, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_11, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_12, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_13, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_14, // @[:@18672.4]
  input  [7:0]  io_inp_data_bits_0_15, // @[:@18672.4]
  input         io_wgt_data_valid, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_0_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_1_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_2_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_3_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_4_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_5_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_6_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_7_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_8_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_9_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_10_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_11_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_12_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_13_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_14_15, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_0, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_1, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_2, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_3, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_4, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_5, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_6, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_7, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_8, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_9, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_10, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_11, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_12, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_13, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_14, // @[:@18672.4]
  input  [7:0]  io_wgt_data_bits_15_15, // @[:@18672.4]
  input         io_acc_i_data_valid, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_0, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_1, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_2, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_3, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_4, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_5, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_6, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_7, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_8, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_9, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_10, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_11, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_12, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_13, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_14, // @[:@18672.4]
  input  [31:0] io_acc_i_data_bits_0_15, // @[:@18672.4]
  output        io_acc_o_data_valid, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_0, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_1, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_2, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_3, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_4, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_5, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_6, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_7, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_8, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_9, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_10, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_11, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_12, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_13, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_14, // @[:@18672.4]
  output [31:0] io_acc_o_data_bits_0_15, // @[:@18672.4]
  output        io_out_data_valid, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_0, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_1, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_2, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_3, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_4, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_5, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_6, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_7, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_8, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_9, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_10, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_11, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_12, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_13, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_14, // @[:@18672.4]
  output [7:0]  io_out_data_bits_0_15 // @[:@18672.4]
);
  wire  dot_0_clock; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_0; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_1; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_2; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_3; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_4; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_5; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_6; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_7; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_8; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_9; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_10; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_11; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_12; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_13; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_14; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_a_15; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_0; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_1; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_2; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_3; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_4; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_5; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_6; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_7; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_8; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_9; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_10; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_11; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_12; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_13; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_14; // @[TensorGemm.scala 153:11:@18674.4]
  wire [7:0] dot_0_io_b_15; // @[TensorGemm.scala 153:11:@18674.4]
  wire [20:0] dot_0_io_y; // @[TensorGemm.scala 153:11:@18674.4]
  wire  dot_1_clock; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_0; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_1; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_2; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_3; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_4; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_5; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_6; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_7; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_8; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_9; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_10; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_11; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_12; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_13; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_14; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_a_15; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_0; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_1; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_2; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_3; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_4; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_5; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_6; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_7; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_8; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_9; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_10; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_11; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_12; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_13; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_14; // @[TensorGemm.scala 153:11:@18677.4]
  wire [7:0] dot_1_io_b_15; // @[TensorGemm.scala 153:11:@18677.4]
  wire [20:0] dot_1_io_y; // @[TensorGemm.scala 153:11:@18677.4]
  wire  dot_2_clock; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_0; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_1; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_2; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_3; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_4; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_5; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_6; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_7; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_8; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_9; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_10; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_11; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_12; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_13; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_14; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_a_15; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_0; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_1; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_2; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_3; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_4; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_5; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_6; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_7; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_8; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_9; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_10; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_11; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_12; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_13; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_14; // @[TensorGemm.scala 153:11:@18680.4]
  wire [7:0] dot_2_io_b_15; // @[TensorGemm.scala 153:11:@18680.4]
  wire [20:0] dot_2_io_y; // @[TensorGemm.scala 153:11:@18680.4]
  wire  dot_3_clock; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_0; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_1; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_2; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_3; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_4; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_5; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_6; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_7; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_8; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_9; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_10; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_11; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_12; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_13; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_14; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_a_15; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_0; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_1; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_2; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_3; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_4; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_5; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_6; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_7; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_8; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_9; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_10; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_11; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_12; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_13; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_14; // @[TensorGemm.scala 153:11:@18683.4]
  wire [7:0] dot_3_io_b_15; // @[TensorGemm.scala 153:11:@18683.4]
  wire [20:0] dot_3_io_y; // @[TensorGemm.scala 153:11:@18683.4]
  wire  dot_4_clock; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_0; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_1; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_2; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_3; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_4; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_5; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_6; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_7; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_8; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_9; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_10; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_11; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_12; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_13; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_14; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_a_15; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_0; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_1; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_2; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_3; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_4; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_5; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_6; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_7; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_8; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_9; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_10; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_11; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_12; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_13; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_14; // @[TensorGemm.scala 153:11:@18686.4]
  wire [7:0] dot_4_io_b_15; // @[TensorGemm.scala 153:11:@18686.4]
  wire [20:0] dot_4_io_y; // @[TensorGemm.scala 153:11:@18686.4]
  wire  dot_5_clock; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_0; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_1; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_2; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_3; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_4; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_5; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_6; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_7; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_8; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_9; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_10; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_11; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_12; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_13; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_14; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_a_15; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_0; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_1; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_2; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_3; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_4; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_5; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_6; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_7; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_8; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_9; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_10; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_11; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_12; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_13; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_14; // @[TensorGemm.scala 153:11:@18689.4]
  wire [7:0] dot_5_io_b_15; // @[TensorGemm.scala 153:11:@18689.4]
  wire [20:0] dot_5_io_y; // @[TensorGemm.scala 153:11:@18689.4]
  wire  dot_6_clock; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_0; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_1; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_2; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_3; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_4; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_5; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_6; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_7; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_8; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_9; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_10; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_11; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_12; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_13; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_14; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_a_15; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_0; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_1; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_2; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_3; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_4; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_5; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_6; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_7; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_8; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_9; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_10; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_11; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_12; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_13; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_14; // @[TensorGemm.scala 153:11:@18692.4]
  wire [7:0] dot_6_io_b_15; // @[TensorGemm.scala 153:11:@18692.4]
  wire [20:0] dot_6_io_y; // @[TensorGemm.scala 153:11:@18692.4]
  wire  dot_7_clock; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_0; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_1; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_2; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_3; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_4; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_5; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_6; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_7; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_8; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_9; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_10; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_11; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_12; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_13; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_14; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_a_15; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_0; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_1; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_2; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_3; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_4; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_5; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_6; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_7; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_8; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_9; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_10; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_11; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_12; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_13; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_14; // @[TensorGemm.scala 153:11:@18695.4]
  wire [7:0] dot_7_io_b_15; // @[TensorGemm.scala 153:11:@18695.4]
  wire [20:0] dot_7_io_y; // @[TensorGemm.scala 153:11:@18695.4]
  wire  dot_8_clock; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_0; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_1; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_2; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_3; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_4; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_5; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_6; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_7; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_8; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_9; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_10; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_11; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_12; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_13; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_14; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_a_15; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_0; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_1; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_2; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_3; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_4; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_5; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_6; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_7; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_8; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_9; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_10; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_11; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_12; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_13; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_14; // @[TensorGemm.scala 153:11:@18698.4]
  wire [7:0] dot_8_io_b_15; // @[TensorGemm.scala 153:11:@18698.4]
  wire [20:0] dot_8_io_y; // @[TensorGemm.scala 153:11:@18698.4]
  wire  dot_9_clock; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_0; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_1; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_2; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_3; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_4; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_5; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_6; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_7; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_8; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_9; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_10; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_11; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_12; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_13; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_14; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_a_15; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_0; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_1; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_2; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_3; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_4; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_5; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_6; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_7; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_8; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_9; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_10; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_11; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_12; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_13; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_14; // @[TensorGemm.scala 153:11:@18701.4]
  wire [7:0] dot_9_io_b_15; // @[TensorGemm.scala 153:11:@18701.4]
  wire [20:0] dot_9_io_y; // @[TensorGemm.scala 153:11:@18701.4]
  wire  dot_10_clock; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_0; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_1; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_2; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_3; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_4; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_5; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_6; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_7; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_8; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_9; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_10; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_11; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_12; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_13; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_14; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_a_15; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_0; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_1; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_2; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_3; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_4; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_5; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_6; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_7; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_8; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_9; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_10; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_11; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_12; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_13; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_14; // @[TensorGemm.scala 153:11:@18704.4]
  wire [7:0] dot_10_io_b_15; // @[TensorGemm.scala 153:11:@18704.4]
  wire [20:0] dot_10_io_y; // @[TensorGemm.scala 153:11:@18704.4]
  wire  dot_11_clock; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_0; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_1; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_2; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_3; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_4; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_5; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_6; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_7; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_8; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_9; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_10; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_11; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_12; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_13; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_14; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_a_15; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_0; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_1; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_2; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_3; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_4; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_5; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_6; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_7; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_8; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_9; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_10; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_11; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_12; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_13; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_14; // @[TensorGemm.scala 153:11:@18707.4]
  wire [7:0] dot_11_io_b_15; // @[TensorGemm.scala 153:11:@18707.4]
  wire [20:0] dot_11_io_y; // @[TensorGemm.scala 153:11:@18707.4]
  wire  dot_12_clock; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_0; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_1; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_2; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_3; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_4; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_5; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_6; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_7; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_8; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_9; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_10; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_11; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_12; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_13; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_14; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_a_15; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_0; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_1; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_2; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_3; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_4; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_5; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_6; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_7; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_8; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_9; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_10; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_11; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_12; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_13; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_14; // @[TensorGemm.scala 153:11:@18710.4]
  wire [7:0] dot_12_io_b_15; // @[TensorGemm.scala 153:11:@18710.4]
  wire [20:0] dot_12_io_y; // @[TensorGemm.scala 153:11:@18710.4]
  wire  dot_13_clock; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_0; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_1; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_2; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_3; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_4; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_5; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_6; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_7; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_8; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_9; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_10; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_11; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_12; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_13; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_14; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_a_15; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_0; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_1; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_2; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_3; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_4; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_5; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_6; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_7; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_8; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_9; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_10; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_11; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_12; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_13; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_14; // @[TensorGemm.scala 153:11:@18713.4]
  wire [7:0] dot_13_io_b_15; // @[TensorGemm.scala 153:11:@18713.4]
  wire [20:0] dot_13_io_y; // @[TensorGemm.scala 153:11:@18713.4]
  wire  dot_14_clock; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_0; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_1; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_2; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_3; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_4; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_5; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_6; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_7; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_8; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_9; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_10; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_11; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_12; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_13; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_14; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_a_15; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_0; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_1; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_2; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_3; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_4; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_5; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_6; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_7; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_8; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_9; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_10; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_11; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_12; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_13; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_14; // @[TensorGemm.scala 153:11:@18716.4]
  wire [7:0] dot_14_io_b_15; // @[TensorGemm.scala 153:11:@18716.4]
  wire [20:0] dot_14_io_y; // @[TensorGemm.scala 153:11:@18716.4]
  wire  dot_15_clock; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_0; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_1; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_2; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_3; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_4; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_5; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_6; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_7; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_8; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_9; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_10; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_11; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_12; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_13; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_14; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_a_15; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_0; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_1; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_2; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_3; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_4; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_5; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_6; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_7; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_8; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_9; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_10; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_11; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_12; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_13; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_14; // @[TensorGemm.scala 153:11:@18719.4]
  wire [7:0] dot_15_io_b_15; // @[TensorGemm.scala 153:11:@18719.4]
  wire [20:0] dot_15_io_y; // @[TensorGemm.scala 153:11:@18719.4]
  wire  acc_0_clock; // @[TensorGemm.scala 156:34:@18722.4]
  wire  acc_0_reset; // @[TensorGemm.scala 156:34:@18722.4]
  wire  acc_0_io_enq_valid; // @[TensorGemm.scala 156:34:@18722.4]
  wire [31:0] acc_0_io_enq_bits; // @[TensorGemm.scala 156:34:@18722.4]
  wire  acc_0_io_deq_valid; // @[TensorGemm.scala 156:34:@18722.4]
  wire [31:0] acc_0_io_deq_bits; // @[TensorGemm.scala 156:34:@18722.4]
  wire  acc_1_clock; // @[TensorGemm.scala 156:34:@18725.4]
  wire  acc_1_reset; // @[TensorGemm.scala 156:34:@18725.4]
  wire  acc_1_io_enq_valid; // @[TensorGemm.scala 156:34:@18725.4]
  wire [31:0] acc_1_io_enq_bits; // @[TensorGemm.scala 156:34:@18725.4]
  wire  acc_1_io_deq_valid; // @[TensorGemm.scala 156:34:@18725.4]
  wire [31:0] acc_1_io_deq_bits; // @[TensorGemm.scala 156:34:@18725.4]
  wire  acc_2_clock; // @[TensorGemm.scala 156:34:@18728.4]
  wire  acc_2_reset; // @[TensorGemm.scala 156:34:@18728.4]
  wire  acc_2_io_enq_valid; // @[TensorGemm.scala 156:34:@18728.4]
  wire [31:0] acc_2_io_enq_bits; // @[TensorGemm.scala 156:34:@18728.4]
  wire  acc_2_io_deq_valid; // @[TensorGemm.scala 156:34:@18728.4]
  wire [31:0] acc_2_io_deq_bits; // @[TensorGemm.scala 156:34:@18728.4]
  wire  acc_3_clock; // @[TensorGemm.scala 156:34:@18731.4]
  wire  acc_3_reset; // @[TensorGemm.scala 156:34:@18731.4]
  wire  acc_3_io_enq_valid; // @[TensorGemm.scala 156:34:@18731.4]
  wire [31:0] acc_3_io_enq_bits; // @[TensorGemm.scala 156:34:@18731.4]
  wire  acc_3_io_deq_valid; // @[TensorGemm.scala 156:34:@18731.4]
  wire [31:0] acc_3_io_deq_bits; // @[TensorGemm.scala 156:34:@18731.4]
  wire  acc_4_clock; // @[TensorGemm.scala 156:34:@18734.4]
  wire  acc_4_reset; // @[TensorGemm.scala 156:34:@18734.4]
  wire  acc_4_io_enq_valid; // @[TensorGemm.scala 156:34:@18734.4]
  wire [31:0] acc_4_io_enq_bits; // @[TensorGemm.scala 156:34:@18734.4]
  wire  acc_4_io_deq_valid; // @[TensorGemm.scala 156:34:@18734.4]
  wire [31:0] acc_4_io_deq_bits; // @[TensorGemm.scala 156:34:@18734.4]
  wire  acc_5_clock; // @[TensorGemm.scala 156:34:@18737.4]
  wire  acc_5_reset; // @[TensorGemm.scala 156:34:@18737.4]
  wire  acc_5_io_enq_valid; // @[TensorGemm.scala 156:34:@18737.4]
  wire [31:0] acc_5_io_enq_bits; // @[TensorGemm.scala 156:34:@18737.4]
  wire  acc_5_io_deq_valid; // @[TensorGemm.scala 156:34:@18737.4]
  wire [31:0] acc_5_io_deq_bits; // @[TensorGemm.scala 156:34:@18737.4]
  wire  acc_6_clock; // @[TensorGemm.scala 156:34:@18740.4]
  wire  acc_6_reset; // @[TensorGemm.scala 156:34:@18740.4]
  wire  acc_6_io_enq_valid; // @[TensorGemm.scala 156:34:@18740.4]
  wire [31:0] acc_6_io_enq_bits; // @[TensorGemm.scala 156:34:@18740.4]
  wire  acc_6_io_deq_valid; // @[TensorGemm.scala 156:34:@18740.4]
  wire [31:0] acc_6_io_deq_bits; // @[TensorGemm.scala 156:34:@18740.4]
  wire  acc_7_clock; // @[TensorGemm.scala 156:34:@18743.4]
  wire  acc_7_reset; // @[TensorGemm.scala 156:34:@18743.4]
  wire  acc_7_io_enq_valid; // @[TensorGemm.scala 156:34:@18743.4]
  wire [31:0] acc_7_io_enq_bits; // @[TensorGemm.scala 156:34:@18743.4]
  wire  acc_7_io_deq_valid; // @[TensorGemm.scala 156:34:@18743.4]
  wire [31:0] acc_7_io_deq_bits; // @[TensorGemm.scala 156:34:@18743.4]
  wire  acc_8_clock; // @[TensorGemm.scala 156:34:@18746.4]
  wire  acc_8_reset; // @[TensorGemm.scala 156:34:@18746.4]
  wire  acc_8_io_enq_valid; // @[TensorGemm.scala 156:34:@18746.4]
  wire [31:0] acc_8_io_enq_bits; // @[TensorGemm.scala 156:34:@18746.4]
  wire  acc_8_io_deq_valid; // @[TensorGemm.scala 156:34:@18746.4]
  wire [31:0] acc_8_io_deq_bits; // @[TensorGemm.scala 156:34:@18746.4]
  wire  acc_9_clock; // @[TensorGemm.scala 156:34:@18749.4]
  wire  acc_9_reset; // @[TensorGemm.scala 156:34:@18749.4]
  wire  acc_9_io_enq_valid; // @[TensorGemm.scala 156:34:@18749.4]
  wire [31:0] acc_9_io_enq_bits; // @[TensorGemm.scala 156:34:@18749.4]
  wire  acc_9_io_deq_valid; // @[TensorGemm.scala 156:34:@18749.4]
  wire [31:0] acc_9_io_deq_bits; // @[TensorGemm.scala 156:34:@18749.4]
  wire  acc_10_clock; // @[TensorGemm.scala 156:34:@18752.4]
  wire  acc_10_reset; // @[TensorGemm.scala 156:34:@18752.4]
  wire  acc_10_io_enq_valid; // @[TensorGemm.scala 156:34:@18752.4]
  wire [31:0] acc_10_io_enq_bits; // @[TensorGemm.scala 156:34:@18752.4]
  wire  acc_10_io_deq_valid; // @[TensorGemm.scala 156:34:@18752.4]
  wire [31:0] acc_10_io_deq_bits; // @[TensorGemm.scala 156:34:@18752.4]
  wire  acc_11_clock; // @[TensorGemm.scala 156:34:@18755.4]
  wire  acc_11_reset; // @[TensorGemm.scala 156:34:@18755.4]
  wire  acc_11_io_enq_valid; // @[TensorGemm.scala 156:34:@18755.4]
  wire [31:0] acc_11_io_enq_bits; // @[TensorGemm.scala 156:34:@18755.4]
  wire  acc_11_io_deq_valid; // @[TensorGemm.scala 156:34:@18755.4]
  wire [31:0] acc_11_io_deq_bits; // @[TensorGemm.scala 156:34:@18755.4]
  wire  acc_12_clock; // @[TensorGemm.scala 156:34:@18758.4]
  wire  acc_12_reset; // @[TensorGemm.scala 156:34:@18758.4]
  wire  acc_12_io_enq_valid; // @[TensorGemm.scala 156:34:@18758.4]
  wire [31:0] acc_12_io_enq_bits; // @[TensorGemm.scala 156:34:@18758.4]
  wire  acc_12_io_deq_valid; // @[TensorGemm.scala 156:34:@18758.4]
  wire [31:0] acc_12_io_deq_bits; // @[TensorGemm.scala 156:34:@18758.4]
  wire  acc_13_clock; // @[TensorGemm.scala 156:34:@18761.4]
  wire  acc_13_reset; // @[TensorGemm.scala 156:34:@18761.4]
  wire  acc_13_io_enq_valid; // @[TensorGemm.scala 156:34:@18761.4]
  wire [31:0] acc_13_io_enq_bits; // @[TensorGemm.scala 156:34:@18761.4]
  wire  acc_13_io_deq_valid; // @[TensorGemm.scala 156:34:@18761.4]
  wire [31:0] acc_13_io_deq_bits; // @[TensorGemm.scala 156:34:@18761.4]
  wire  acc_14_clock; // @[TensorGemm.scala 156:34:@18764.4]
  wire  acc_14_reset; // @[TensorGemm.scala 156:34:@18764.4]
  wire  acc_14_io_enq_valid; // @[TensorGemm.scala 156:34:@18764.4]
  wire [31:0] acc_14_io_enq_bits; // @[TensorGemm.scala 156:34:@18764.4]
  wire  acc_14_io_deq_valid; // @[TensorGemm.scala 156:34:@18764.4]
  wire [31:0] acc_14_io_deq_bits; // @[TensorGemm.scala 156:34:@18764.4]
  wire  acc_15_clock; // @[TensorGemm.scala 156:34:@18767.4]
  wire  acc_15_reset; // @[TensorGemm.scala 156:34:@18767.4]
  wire  acc_15_io_enq_valid; // @[TensorGemm.scala 156:34:@18767.4]
  wire [31:0] acc_15_io_enq_bits; // @[TensorGemm.scala 156:34:@18767.4]
  wire  acc_15_io_deq_valid; // @[TensorGemm.scala 156:34:@18767.4]
  wire [31:0] acc_15_io_deq_bits; // @[TensorGemm.scala 156:34:@18767.4]
  wire  _T_6016; // @[TensorGemm.scala 161:46:@18787.4]
  wire  _T_6017; // @[TensorGemm.scala 161:66:@18788.4]
  wire  _T_6018; // @[TensorGemm.scala 161:90:@18789.4]
  wire [31:0] _T_6052; // @[TensorGemm.scala 167:34:@18857.4]
  wire [31:0] _GEN_0; // @[TensorGemm.scala 167:41:@18858.4]
  wire [32:0] _T_6053; // @[TensorGemm.scala 167:41:@18858.4]
  wire [31:0] _T_6054; // @[TensorGemm.scala 167:41:@18859.4]
  wire [31:0] add_0; // @[TensorGemm.scala 167:41:@18860.4]
  wire [31:0] _T_6057; // @[TensorGemm.scala 168:59:@18862.4]
  wire [31:0] _T_6096; // @[TensorGemm.scala 167:34:@18938.4]
  wire [31:0] _GEN_1; // @[TensorGemm.scala 167:41:@18939.4]
  wire [32:0] _T_6097; // @[TensorGemm.scala 167:41:@18939.4]
  wire [31:0] _T_6098; // @[TensorGemm.scala 167:41:@18940.4]
  wire [31:0] add_1; // @[TensorGemm.scala 167:41:@18941.4]
  wire [31:0] _T_6101; // @[TensorGemm.scala 168:59:@18943.4]
  wire [31:0] _T_6140; // @[TensorGemm.scala 167:34:@19019.4]
  wire [31:0] _GEN_2; // @[TensorGemm.scala 167:41:@19020.4]
  wire [32:0] _T_6141; // @[TensorGemm.scala 167:41:@19020.4]
  wire [31:0] _T_6142; // @[TensorGemm.scala 167:41:@19021.4]
  wire [31:0] add_2; // @[TensorGemm.scala 167:41:@19022.4]
  wire [31:0] _T_6145; // @[TensorGemm.scala 168:59:@19024.4]
  wire [31:0] _T_6184; // @[TensorGemm.scala 167:34:@19100.4]
  wire [31:0] _GEN_3; // @[TensorGemm.scala 167:41:@19101.4]
  wire [32:0] _T_6185; // @[TensorGemm.scala 167:41:@19101.4]
  wire [31:0] _T_6186; // @[TensorGemm.scala 167:41:@19102.4]
  wire [31:0] add_3; // @[TensorGemm.scala 167:41:@19103.4]
  wire [31:0] _T_6189; // @[TensorGemm.scala 168:59:@19105.4]
  wire [31:0] _T_6228; // @[TensorGemm.scala 167:34:@19181.4]
  wire [31:0] _GEN_4; // @[TensorGemm.scala 167:41:@19182.4]
  wire [32:0] _T_6229; // @[TensorGemm.scala 167:41:@19182.4]
  wire [31:0] _T_6230; // @[TensorGemm.scala 167:41:@19183.4]
  wire [31:0] add_4; // @[TensorGemm.scala 167:41:@19184.4]
  wire [31:0] _T_6233; // @[TensorGemm.scala 168:59:@19186.4]
  wire [31:0] _T_6272; // @[TensorGemm.scala 167:34:@19262.4]
  wire [31:0] _GEN_5; // @[TensorGemm.scala 167:41:@19263.4]
  wire [32:0] _T_6273; // @[TensorGemm.scala 167:41:@19263.4]
  wire [31:0] _T_6274; // @[TensorGemm.scala 167:41:@19264.4]
  wire [31:0] add_5; // @[TensorGemm.scala 167:41:@19265.4]
  wire [31:0] _T_6277; // @[TensorGemm.scala 168:59:@19267.4]
  wire [31:0] _T_6316; // @[TensorGemm.scala 167:34:@19343.4]
  wire [31:0] _GEN_6; // @[TensorGemm.scala 167:41:@19344.4]
  wire [32:0] _T_6317; // @[TensorGemm.scala 167:41:@19344.4]
  wire [31:0] _T_6318; // @[TensorGemm.scala 167:41:@19345.4]
  wire [31:0] add_6; // @[TensorGemm.scala 167:41:@19346.4]
  wire [31:0] _T_6321; // @[TensorGemm.scala 168:59:@19348.4]
  wire [31:0] _T_6360; // @[TensorGemm.scala 167:34:@19424.4]
  wire [31:0] _GEN_7; // @[TensorGemm.scala 167:41:@19425.4]
  wire [32:0] _T_6361; // @[TensorGemm.scala 167:41:@19425.4]
  wire [31:0] _T_6362; // @[TensorGemm.scala 167:41:@19426.4]
  wire [31:0] add_7; // @[TensorGemm.scala 167:41:@19427.4]
  wire [31:0] _T_6365; // @[TensorGemm.scala 168:59:@19429.4]
  wire [31:0] _T_6404; // @[TensorGemm.scala 167:34:@19505.4]
  wire [31:0] _GEN_8; // @[TensorGemm.scala 167:41:@19506.4]
  wire [32:0] _T_6405; // @[TensorGemm.scala 167:41:@19506.4]
  wire [31:0] _T_6406; // @[TensorGemm.scala 167:41:@19507.4]
  wire [31:0] add_8; // @[TensorGemm.scala 167:41:@19508.4]
  wire [31:0] _T_6409; // @[TensorGemm.scala 168:59:@19510.4]
  wire [31:0] _T_6448; // @[TensorGemm.scala 167:34:@19586.4]
  wire [31:0] _GEN_9; // @[TensorGemm.scala 167:41:@19587.4]
  wire [32:0] _T_6449; // @[TensorGemm.scala 167:41:@19587.4]
  wire [31:0] _T_6450; // @[TensorGemm.scala 167:41:@19588.4]
  wire [31:0] add_9; // @[TensorGemm.scala 167:41:@19589.4]
  wire [31:0] _T_6453; // @[TensorGemm.scala 168:59:@19591.4]
  wire [31:0] _T_6492; // @[TensorGemm.scala 167:34:@19667.4]
  wire [31:0] _GEN_10; // @[TensorGemm.scala 167:41:@19668.4]
  wire [32:0] _T_6493; // @[TensorGemm.scala 167:41:@19668.4]
  wire [31:0] _T_6494; // @[TensorGemm.scala 167:41:@19669.4]
  wire [31:0] add_10; // @[TensorGemm.scala 167:41:@19670.4]
  wire [31:0] _T_6497; // @[TensorGemm.scala 168:59:@19672.4]
  wire [31:0] _T_6536; // @[TensorGemm.scala 167:34:@19748.4]
  wire [31:0] _GEN_11; // @[TensorGemm.scala 167:41:@19749.4]
  wire [32:0] _T_6537; // @[TensorGemm.scala 167:41:@19749.4]
  wire [31:0] _T_6538; // @[TensorGemm.scala 167:41:@19750.4]
  wire [31:0] add_11; // @[TensorGemm.scala 167:41:@19751.4]
  wire [31:0] _T_6541; // @[TensorGemm.scala 168:59:@19753.4]
  wire [31:0] _T_6580; // @[TensorGemm.scala 167:34:@19829.4]
  wire [31:0] _GEN_12; // @[TensorGemm.scala 167:41:@19830.4]
  wire [32:0] _T_6581; // @[TensorGemm.scala 167:41:@19830.4]
  wire [31:0] _T_6582; // @[TensorGemm.scala 167:41:@19831.4]
  wire [31:0] add_12; // @[TensorGemm.scala 167:41:@19832.4]
  wire [31:0] _T_6585; // @[TensorGemm.scala 168:59:@19834.4]
  wire [31:0] _T_6624; // @[TensorGemm.scala 167:34:@19910.4]
  wire [31:0] _GEN_13; // @[TensorGemm.scala 167:41:@19911.4]
  wire [32:0] _T_6625; // @[TensorGemm.scala 167:41:@19911.4]
  wire [31:0] _T_6626; // @[TensorGemm.scala 167:41:@19912.4]
  wire [31:0] add_13; // @[TensorGemm.scala 167:41:@19913.4]
  wire [31:0] _T_6629; // @[TensorGemm.scala 168:59:@19915.4]
  wire [31:0] _T_6668; // @[TensorGemm.scala 167:34:@19991.4]
  wire [31:0] _GEN_14; // @[TensorGemm.scala 167:41:@19992.4]
  wire [32:0] _T_6669; // @[TensorGemm.scala 167:41:@19992.4]
  wire [31:0] _T_6670; // @[TensorGemm.scala 167:41:@19993.4]
  wire [31:0] add_14; // @[TensorGemm.scala 167:41:@19994.4]
  wire [31:0] _T_6673; // @[TensorGemm.scala 168:59:@19996.4]
  wire [31:0] _T_6712; // @[TensorGemm.scala 167:34:@20072.4]
  wire [31:0] _GEN_15; // @[TensorGemm.scala 167:41:@20073.4]
  wire [32:0] _T_6713; // @[TensorGemm.scala 167:41:@20073.4]
  wire [31:0] _T_6714; // @[TensorGemm.scala 167:41:@20074.4]
  wire [31:0] add_15; // @[TensorGemm.scala 167:41:@20075.4]
  wire [31:0] _T_6717; // @[TensorGemm.scala 168:59:@20077.4]
  wire  vld_1; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@18948.4]
  wire  vld_0; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@18867.4]
  wire  vld_3; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19110.4]
  wire  vld_2; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19029.4]
  wire  vld_5; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19272.4]
  wire  vld_4; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19191.4]
  wire  vld_7; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19434.4]
  wire  vld_6; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19353.4]
  wire [7:0] _T_6726; // @[TensorGemm.scala 172:30:@20089.4]
  wire  vld_9; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19596.4]
  wire  vld_8; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19515.4]
  wire  vld_11; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19758.4]
  wire  vld_10; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19677.4]
  wire  vld_13; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19920.4]
  wire  vld_12; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19839.4]
  wire  vld_15; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@20082.4]
  wire  vld_14; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@20001.4]
  wire [15:0] _T_6734; // @[TensorGemm.scala 172:30:@20097.4]
  wire [15:0] _T_6735; // @[TensorGemm.scala 172:37:@20098.4]
  wire  _T_6737; // @[TensorGemm.scala 172:37:@20099.4]
  DotProduct dot_0 ( // @[TensorGemm.scala 153:11:@18674.4]
    .clock(dot_0_clock),
    .io_a_0(dot_0_io_a_0),
    .io_a_1(dot_0_io_a_1),
    .io_a_2(dot_0_io_a_2),
    .io_a_3(dot_0_io_a_3),
    .io_a_4(dot_0_io_a_4),
    .io_a_5(dot_0_io_a_5),
    .io_a_6(dot_0_io_a_6),
    .io_a_7(dot_0_io_a_7),
    .io_a_8(dot_0_io_a_8),
    .io_a_9(dot_0_io_a_9),
    .io_a_10(dot_0_io_a_10),
    .io_a_11(dot_0_io_a_11),
    .io_a_12(dot_0_io_a_12),
    .io_a_13(dot_0_io_a_13),
    .io_a_14(dot_0_io_a_14),
    .io_a_15(dot_0_io_a_15),
    .io_b_0(dot_0_io_b_0),
    .io_b_1(dot_0_io_b_1),
    .io_b_2(dot_0_io_b_2),
    .io_b_3(dot_0_io_b_3),
    .io_b_4(dot_0_io_b_4),
    .io_b_5(dot_0_io_b_5),
    .io_b_6(dot_0_io_b_6),
    .io_b_7(dot_0_io_b_7),
    .io_b_8(dot_0_io_b_8),
    .io_b_9(dot_0_io_b_9),
    .io_b_10(dot_0_io_b_10),
    .io_b_11(dot_0_io_b_11),
    .io_b_12(dot_0_io_b_12),
    .io_b_13(dot_0_io_b_13),
    .io_b_14(dot_0_io_b_14),
    .io_b_15(dot_0_io_b_15),
    .io_y(dot_0_io_y)
  );
  DotProduct dot_1 ( // @[TensorGemm.scala 153:11:@18677.4]
    .clock(dot_1_clock),
    .io_a_0(dot_1_io_a_0),
    .io_a_1(dot_1_io_a_1),
    .io_a_2(dot_1_io_a_2),
    .io_a_3(dot_1_io_a_3),
    .io_a_4(dot_1_io_a_4),
    .io_a_5(dot_1_io_a_5),
    .io_a_6(dot_1_io_a_6),
    .io_a_7(dot_1_io_a_7),
    .io_a_8(dot_1_io_a_8),
    .io_a_9(dot_1_io_a_9),
    .io_a_10(dot_1_io_a_10),
    .io_a_11(dot_1_io_a_11),
    .io_a_12(dot_1_io_a_12),
    .io_a_13(dot_1_io_a_13),
    .io_a_14(dot_1_io_a_14),
    .io_a_15(dot_1_io_a_15),
    .io_b_0(dot_1_io_b_0),
    .io_b_1(dot_1_io_b_1),
    .io_b_2(dot_1_io_b_2),
    .io_b_3(dot_1_io_b_3),
    .io_b_4(dot_1_io_b_4),
    .io_b_5(dot_1_io_b_5),
    .io_b_6(dot_1_io_b_6),
    .io_b_7(dot_1_io_b_7),
    .io_b_8(dot_1_io_b_8),
    .io_b_9(dot_1_io_b_9),
    .io_b_10(dot_1_io_b_10),
    .io_b_11(dot_1_io_b_11),
    .io_b_12(dot_1_io_b_12),
    .io_b_13(dot_1_io_b_13),
    .io_b_14(dot_1_io_b_14),
    .io_b_15(dot_1_io_b_15),
    .io_y(dot_1_io_y)
  );
  DotProduct dot_2 ( // @[TensorGemm.scala 153:11:@18680.4]
    .clock(dot_2_clock),
    .io_a_0(dot_2_io_a_0),
    .io_a_1(dot_2_io_a_1),
    .io_a_2(dot_2_io_a_2),
    .io_a_3(dot_2_io_a_3),
    .io_a_4(dot_2_io_a_4),
    .io_a_5(dot_2_io_a_5),
    .io_a_6(dot_2_io_a_6),
    .io_a_7(dot_2_io_a_7),
    .io_a_8(dot_2_io_a_8),
    .io_a_9(dot_2_io_a_9),
    .io_a_10(dot_2_io_a_10),
    .io_a_11(dot_2_io_a_11),
    .io_a_12(dot_2_io_a_12),
    .io_a_13(dot_2_io_a_13),
    .io_a_14(dot_2_io_a_14),
    .io_a_15(dot_2_io_a_15),
    .io_b_0(dot_2_io_b_0),
    .io_b_1(dot_2_io_b_1),
    .io_b_2(dot_2_io_b_2),
    .io_b_3(dot_2_io_b_3),
    .io_b_4(dot_2_io_b_4),
    .io_b_5(dot_2_io_b_5),
    .io_b_6(dot_2_io_b_6),
    .io_b_7(dot_2_io_b_7),
    .io_b_8(dot_2_io_b_8),
    .io_b_9(dot_2_io_b_9),
    .io_b_10(dot_2_io_b_10),
    .io_b_11(dot_2_io_b_11),
    .io_b_12(dot_2_io_b_12),
    .io_b_13(dot_2_io_b_13),
    .io_b_14(dot_2_io_b_14),
    .io_b_15(dot_2_io_b_15),
    .io_y(dot_2_io_y)
  );
  DotProduct dot_3 ( // @[TensorGemm.scala 153:11:@18683.4]
    .clock(dot_3_clock),
    .io_a_0(dot_3_io_a_0),
    .io_a_1(dot_3_io_a_1),
    .io_a_2(dot_3_io_a_2),
    .io_a_3(dot_3_io_a_3),
    .io_a_4(dot_3_io_a_4),
    .io_a_5(dot_3_io_a_5),
    .io_a_6(dot_3_io_a_6),
    .io_a_7(dot_3_io_a_7),
    .io_a_8(dot_3_io_a_8),
    .io_a_9(dot_3_io_a_9),
    .io_a_10(dot_3_io_a_10),
    .io_a_11(dot_3_io_a_11),
    .io_a_12(dot_3_io_a_12),
    .io_a_13(dot_3_io_a_13),
    .io_a_14(dot_3_io_a_14),
    .io_a_15(dot_3_io_a_15),
    .io_b_0(dot_3_io_b_0),
    .io_b_1(dot_3_io_b_1),
    .io_b_2(dot_3_io_b_2),
    .io_b_3(dot_3_io_b_3),
    .io_b_4(dot_3_io_b_4),
    .io_b_5(dot_3_io_b_5),
    .io_b_6(dot_3_io_b_6),
    .io_b_7(dot_3_io_b_7),
    .io_b_8(dot_3_io_b_8),
    .io_b_9(dot_3_io_b_9),
    .io_b_10(dot_3_io_b_10),
    .io_b_11(dot_3_io_b_11),
    .io_b_12(dot_3_io_b_12),
    .io_b_13(dot_3_io_b_13),
    .io_b_14(dot_3_io_b_14),
    .io_b_15(dot_3_io_b_15),
    .io_y(dot_3_io_y)
  );
  DotProduct dot_4 ( // @[TensorGemm.scala 153:11:@18686.4]
    .clock(dot_4_clock),
    .io_a_0(dot_4_io_a_0),
    .io_a_1(dot_4_io_a_1),
    .io_a_2(dot_4_io_a_2),
    .io_a_3(dot_4_io_a_3),
    .io_a_4(dot_4_io_a_4),
    .io_a_5(dot_4_io_a_5),
    .io_a_6(dot_4_io_a_6),
    .io_a_7(dot_4_io_a_7),
    .io_a_8(dot_4_io_a_8),
    .io_a_9(dot_4_io_a_9),
    .io_a_10(dot_4_io_a_10),
    .io_a_11(dot_4_io_a_11),
    .io_a_12(dot_4_io_a_12),
    .io_a_13(dot_4_io_a_13),
    .io_a_14(dot_4_io_a_14),
    .io_a_15(dot_4_io_a_15),
    .io_b_0(dot_4_io_b_0),
    .io_b_1(dot_4_io_b_1),
    .io_b_2(dot_4_io_b_2),
    .io_b_3(dot_4_io_b_3),
    .io_b_4(dot_4_io_b_4),
    .io_b_5(dot_4_io_b_5),
    .io_b_6(dot_4_io_b_6),
    .io_b_7(dot_4_io_b_7),
    .io_b_8(dot_4_io_b_8),
    .io_b_9(dot_4_io_b_9),
    .io_b_10(dot_4_io_b_10),
    .io_b_11(dot_4_io_b_11),
    .io_b_12(dot_4_io_b_12),
    .io_b_13(dot_4_io_b_13),
    .io_b_14(dot_4_io_b_14),
    .io_b_15(dot_4_io_b_15),
    .io_y(dot_4_io_y)
  );
  DotProduct dot_5 ( // @[TensorGemm.scala 153:11:@18689.4]
    .clock(dot_5_clock),
    .io_a_0(dot_5_io_a_0),
    .io_a_1(dot_5_io_a_1),
    .io_a_2(dot_5_io_a_2),
    .io_a_3(dot_5_io_a_3),
    .io_a_4(dot_5_io_a_4),
    .io_a_5(dot_5_io_a_5),
    .io_a_6(dot_5_io_a_6),
    .io_a_7(dot_5_io_a_7),
    .io_a_8(dot_5_io_a_8),
    .io_a_9(dot_5_io_a_9),
    .io_a_10(dot_5_io_a_10),
    .io_a_11(dot_5_io_a_11),
    .io_a_12(dot_5_io_a_12),
    .io_a_13(dot_5_io_a_13),
    .io_a_14(dot_5_io_a_14),
    .io_a_15(dot_5_io_a_15),
    .io_b_0(dot_5_io_b_0),
    .io_b_1(dot_5_io_b_1),
    .io_b_2(dot_5_io_b_2),
    .io_b_3(dot_5_io_b_3),
    .io_b_4(dot_5_io_b_4),
    .io_b_5(dot_5_io_b_5),
    .io_b_6(dot_5_io_b_6),
    .io_b_7(dot_5_io_b_7),
    .io_b_8(dot_5_io_b_8),
    .io_b_9(dot_5_io_b_9),
    .io_b_10(dot_5_io_b_10),
    .io_b_11(dot_5_io_b_11),
    .io_b_12(dot_5_io_b_12),
    .io_b_13(dot_5_io_b_13),
    .io_b_14(dot_5_io_b_14),
    .io_b_15(dot_5_io_b_15),
    .io_y(dot_5_io_y)
  );
  DotProduct dot_6 ( // @[TensorGemm.scala 153:11:@18692.4]
    .clock(dot_6_clock),
    .io_a_0(dot_6_io_a_0),
    .io_a_1(dot_6_io_a_1),
    .io_a_2(dot_6_io_a_2),
    .io_a_3(dot_6_io_a_3),
    .io_a_4(dot_6_io_a_4),
    .io_a_5(dot_6_io_a_5),
    .io_a_6(dot_6_io_a_6),
    .io_a_7(dot_6_io_a_7),
    .io_a_8(dot_6_io_a_8),
    .io_a_9(dot_6_io_a_9),
    .io_a_10(dot_6_io_a_10),
    .io_a_11(dot_6_io_a_11),
    .io_a_12(dot_6_io_a_12),
    .io_a_13(dot_6_io_a_13),
    .io_a_14(dot_6_io_a_14),
    .io_a_15(dot_6_io_a_15),
    .io_b_0(dot_6_io_b_0),
    .io_b_1(dot_6_io_b_1),
    .io_b_2(dot_6_io_b_2),
    .io_b_3(dot_6_io_b_3),
    .io_b_4(dot_6_io_b_4),
    .io_b_5(dot_6_io_b_5),
    .io_b_6(dot_6_io_b_6),
    .io_b_7(dot_6_io_b_7),
    .io_b_8(dot_6_io_b_8),
    .io_b_9(dot_6_io_b_9),
    .io_b_10(dot_6_io_b_10),
    .io_b_11(dot_6_io_b_11),
    .io_b_12(dot_6_io_b_12),
    .io_b_13(dot_6_io_b_13),
    .io_b_14(dot_6_io_b_14),
    .io_b_15(dot_6_io_b_15),
    .io_y(dot_6_io_y)
  );
  DotProduct dot_7 ( // @[TensorGemm.scala 153:11:@18695.4]
    .clock(dot_7_clock),
    .io_a_0(dot_7_io_a_0),
    .io_a_1(dot_7_io_a_1),
    .io_a_2(dot_7_io_a_2),
    .io_a_3(dot_7_io_a_3),
    .io_a_4(dot_7_io_a_4),
    .io_a_5(dot_7_io_a_5),
    .io_a_6(dot_7_io_a_6),
    .io_a_7(dot_7_io_a_7),
    .io_a_8(dot_7_io_a_8),
    .io_a_9(dot_7_io_a_9),
    .io_a_10(dot_7_io_a_10),
    .io_a_11(dot_7_io_a_11),
    .io_a_12(dot_7_io_a_12),
    .io_a_13(dot_7_io_a_13),
    .io_a_14(dot_7_io_a_14),
    .io_a_15(dot_7_io_a_15),
    .io_b_0(dot_7_io_b_0),
    .io_b_1(dot_7_io_b_1),
    .io_b_2(dot_7_io_b_2),
    .io_b_3(dot_7_io_b_3),
    .io_b_4(dot_7_io_b_4),
    .io_b_5(dot_7_io_b_5),
    .io_b_6(dot_7_io_b_6),
    .io_b_7(dot_7_io_b_7),
    .io_b_8(dot_7_io_b_8),
    .io_b_9(dot_7_io_b_9),
    .io_b_10(dot_7_io_b_10),
    .io_b_11(dot_7_io_b_11),
    .io_b_12(dot_7_io_b_12),
    .io_b_13(dot_7_io_b_13),
    .io_b_14(dot_7_io_b_14),
    .io_b_15(dot_7_io_b_15),
    .io_y(dot_7_io_y)
  );
  DotProduct dot_8 ( // @[TensorGemm.scala 153:11:@18698.4]
    .clock(dot_8_clock),
    .io_a_0(dot_8_io_a_0),
    .io_a_1(dot_8_io_a_1),
    .io_a_2(dot_8_io_a_2),
    .io_a_3(dot_8_io_a_3),
    .io_a_4(dot_8_io_a_4),
    .io_a_5(dot_8_io_a_5),
    .io_a_6(dot_8_io_a_6),
    .io_a_7(dot_8_io_a_7),
    .io_a_8(dot_8_io_a_8),
    .io_a_9(dot_8_io_a_9),
    .io_a_10(dot_8_io_a_10),
    .io_a_11(dot_8_io_a_11),
    .io_a_12(dot_8_io_a_12),
    .io_a_13(dot_8_io_a_13),
    .io_a_14(dot_8_io_a_14),
    .io_a_15(dot_8_io_a_15),
    .io_b_0(dot_8_io_b_0),
    .io_b_1(dot_8_io_b_1),
    .io_b_2(dot_8_io_b_2),
    .io_b_3(dot_8_io_b_3),
    .io_b_4(dot_8_io_b_4),
    .io_b_5(dot_8_io_b_5),
    .io_b_6(dot_8_io_b_6),
    .io_b_7(dot_8_io_b_7),
    .io_b_8(dot_8_io_b_8),
    .io_b_9(dot_8_io_b_9),
    .io_b_10(dot_8_io_b_10),
    .io_b_11(dot_8_io_b_11),
    .io_b_12(dot_8_io_b_12),
    .io_b_13(dot_8_io_b_13),
    .io_b_14(dot_8_io_b_14),
    .io_b_15(dot_8_io_b_15),
    .io_y(dot_8_io_y)
  );
  DotProduct dot_9 ( // @[TensorGemm.scala 153:11:@18701.4]
    .clock(dot_9_clock),
    .io_a_0(dot_9_io_a_0),
    .io_a_1(dot_9_io_a_1),
    .io_a_2(dot_9_io_a_2),
    .io_a_3(dot_9_io_a_3),
    .io_a_4(dot_9_io_a_4),
    .io_a_5(dot_9_io_a_5),
    .io_a_6(dot_9_io_a_6),
    .io_a_7(dot_9_io_a_7),
    .io_a_8(dot_9_io_a_8),
    .io_a_9(dot_9_io_a_9),
    .io_a_10(dot_9_io_a_10),
    .io_a_11(dot_9_io_a_11),
    .io_a_12(dot_9_io_a_12),
    .io_a_13(dot_9_io_a_13),
    .io_a_14(dot_9_io_a_14),
    .io_a_15(dot_9_io_a_15),
    .io_b_0(dot_9_io_b_0),
    .io_b_1(dot_9_io_b_1),
    .io_b_2(dot_9_io_b_2),
    .io_b_3(dot_9_io_b_3),
    .io_b_4(dot_9_io_b_4),
    .io_b_5(dot_9_io_b_5),
    .io_b_6(dot_9_io_b_6),
    .io_b_7(dot_9_io_b_7),
    .io_b_8(dot_9_io_b_8),
    .io_b_9(dot_9_io_b_9),
    .io_b_10(dot_9_io_b_10),
    .io_b_11(dot_9_io_b_11),
    .io_b_12(dot_9_io_b_12),
    .io_b_13(dot_9_io_b_13),
    .io_b_14(dot_9_io_b_14),
    .io_b_15(dot_9_io_b_15),
    .io_y(dot_9_io_y)
  );
  DotProduct dot_10 ( // @[TensorGemm.scala 153:11:@18704.4]
    .clock(dot_10_clock),
    .io_a_0(dot_10_io_a_0),
    .io_a_1(dot_10_io_a_1),
    .io_a_2(dot_10_io_a_2),
    .io_a_3(dot_10_io_a_3),
    .io_a_4(dot_10_io_a_4),
    .io_a_5(dot_10_io_a_5),
    .io_a_6(dot_10_io_a_6),
    .io_a_7(dot_10_io_a_7),
    .io_a_8(dot_10_io_a_8),
    .io_a_9(dot_10_io_a_9),
    .io_a_10(dot_10_io_a_10),
    .io_a_11(dot_10_io_a_11),
    .io_a_12(dot_10_io_a_12),
    .io_a_13(dot_10_io_a_13),
    .io_a_14(dot_10_io_a_14),
    .io_a_15(dot_10_io_a_15),
    .io_b_0(dot_10_io_b_0),
    .io_b_1(dot_10_io_b_1),
    .io_b_2(dot_10_io_b_2),
    .io_b_3(dot_10_io_b_3),
    .io_b_4(dot_10_io_b_4),
    .io_b_5(dot_10_io_b_5),
    .io_b_6(dot_10_io_b_6),
    .io_b_7(dot_10_io_b_7),
    .io_b_8(dot_10_io_b_8),
    .io_b_9(dot_10_io_b_9),
    .io_b_10(dot_10_io_b_10),
    .io_b_11(dot_10_io_b_11),
    .io_b_12(dot_10_io_b_12),
    .io_b_13(dot_10_io_b_13),
    .io_b_14(dot_10_io_b_14),
    .io_b_15(dot_10_io_b_15),
    .io_y(dot_10_io_y)
  );
  DotProduct dot_11 ( // @[TensorGemm.scala 153:11:@18707.4]
    .clock(dot_11_clock),
    .io_a_0(dot_11_io_a_0),
    .io_a_1(dot_11_io_a_1),
    .io_a_2(dot_11_io_a_2),
    .io_a_3(dot_11_io_a_3),
    .io_a_4(dot_11_io_a_4),
    .io_a_5(dot_11_io_a_5),
    .io_a_6(dot_11_io_a_6),
    .io_a_7(dot_11_io_a_7),
    .io_a_8(dot_11_io_a_8),
    .io_a_9(dot_11_io_a_9),
    .io_a_10(dot_11_io_a_10),
    .io_a_11(dot_11_io_a_11),
    .io_a_12(dot_11_io_a_12),
    .io_a_13(dot_11_io_a_13),
    .io_a_14(dot_11_io_a_14),
    .io_a_15(dot_11_io_a_15),
    .io_b_0(dot_11_io_b_0),
    .io_b_1(dot_11_io_b_1),
    .io_b_2(dot_11_io_b_2),
    .io_b_3(dot_11_io_b_3),
    .io_b_4(dot_11_io_b_4),
    .io_b_5(dot_11_io_b_5),
    .io_b_6(dot_11_io_b_6),
    .io_b_7(dot_11_io_b_7),
    .io_b_8(dot_11_io_b_8),
    .io_b_9(dot_11_io_b_9),
    .io_b_10(dot_11_io_b_10),
    .io_b_11(dot_11_io_b_11),
    .io_b_12(dot_11_io_b_12),
    .io_b_13(dot_11_io_b_13),
    .io_b_14(dot_11_io_b_14),
    .io_b_15(dot_11_io_b_15),
    .io_y(dot_11_io_y)
  );
  DotProduct dot_12 ( // @[TensorGemm.scala 153:11:@18710.4]
    .clock(dot_12_clock),
    .io_a_0(dot_12_io_a_0),
    .io_a_1(dot_12_io_a_1),
    .io_a_2(dot_12_io_a_2),
    .io_a_3(dot_12_io_a_3),
    .io_a_4(dot_12_io_a_4),
    .io_a_5(dot_12_io_a_5),
    .io_a_6(dot_12_io_a_6),
    .io_a_7(dot_12_io_a_7),
    .io_a_8(dot_12_io_a_8),
    .io_a_9(dot_12_io_a_9),
    .io_a_10(dot_12_io_a_10),
    .io_a_11(dot_12_io_a_11),
    .io_a_12(dot_12_io_a_12),
    .io_a_13(dot_12_io_a_13),
    .io_a_14(dot_12_io_a_14),
    .io_a_15(dot_12_io_a_15),
    .io_b_0(dot_12_io_b_0),
    .io_b_1(dot_12_io_b_1),
    .io_b_2(dot_12_io_b_2),
    .io_b_3(dot_12_io_b_3),
    .io_b_4(dot_12_io_b_4),
    .io_b_5(dot_12_io_b_5),
    .io_b_6(dot_12_io_b_6),
    .io_b_7(dot_12_io_b_7),
    .io_b_8(dot_12_io_b_8),
    .io_b_9(dot_12_io_b_9),
    .io_b_10(dot_12_io_b_10),
    .io_b_11(dot_12_io_b_11),
    .io_b_12(dot_12_io_b_12),
    .io_b_13(dot_12_io_b_13),
    .io_b_14(dot_12_io_b_14),
    .io_b_15(dot_12_io_b_15),
    .io_y(dot_12_io_y)
  );
  DotProduct dot_13 ( // @[TensorGemm.scala 153:11:@18713.4]
    .clock(dot_13_clock),
    .io_a_0(dot_13_io_a_0),
    .io_a_1(dot_13_io_a_1),
    .io_a_2(dot_13_io_a_2),
    .io_a_3(dot_13_io_a_3),
    .io_a_4(dot_13_io_a_4),
    .io_a_5(dot_13_io_a_5),
    .io_a_6(dot_13_io_a_6),
    .io_a_7(dot_13_io_a_7),
    .io_a_8(dot_13_io_a_8),
    .io_a_9(dot_13_io_a_9),
    .io_a_10(dot_13_io_a_10),
    .io_a_11(dot_13_io_a_11),
    .io_a_12(dot_13_io_a_12),
    .io_a_13(dot_13_io_a_13),
    .io_a_14(dot_13_io_a_14),
    .io_a_15(dot_13_io_a_15),
    .io_b_0(dot_13_io_b_0),
    .io_b_1(dot_13_io_b_1),
    .io_b_2(dot_13_io_b_2),
    .io_b_3(dot_13_io_b_3),
    .io_b_4(dot_13_io_b_4),
    .io_b_5(dot_13_io_b_5),
    .io_b_6(dot_13_io_b_6),
    .io_b_7(dot_13_io_b_7),
    .io_b_8(dot_13_io_b_8),
    .io_b_9(dot_13_io_b_9),
    .io_b_10(dot_13_io_b_10),
    .io_b_11(dot_13_io_b_11),
    .io_b_12(dot_13_io_b_12),
    .io_b_13(dot_13_io_b_13),
    .io_b_14(dot_13_io_b_14),
    .io_b_15(dot_13_io_b_15),
    .io_y(dot_13_io_y)
  );
  DotProduct dot_14 ( // @[TensorGemm.scala 153:11:@18716.4]
    .clock(dot_14_clock),
    .io_a_0(dot_14_io_a_0),
    .io_a_1(dot_14_io_a_1),
    .io_a_2(dot_14_io_a_2),
    .io_a_3(dot_14_io_a_3),
    .io_a_4(dot_14_io_a_4),
    .io_a_5(dot_14_io_a_5),
    .io_a_6(dot_14_io_a_6),
    .io_a_7(dot_14_io_a_7),
    .io_a_8(dot_14_io_a_8),
    .io_a_9(dot_14_io_a_9),
    .io_a_10(dot_14_io_a_10),
    .io_a_11(dot_14_io_a_11),
    .io_a_12(dot_14_io_a_12),
    .io_a_13(dot_14_io_a_13),
    .io_a_14(dot_14_io_a_14),
    .io_a_15(dot_14_io_a_15),
    .io_b_0(dot_14_io_b_0),
    .io_b_1(dot_14_io_b_1),
    .io_b_2(dot_14_io_b_2),
    .io_b_3(dot_14_io_b_3),
    .io_b_4(dot_14_io_b_4),
    .io_b_5(dot_14_io_b_5),
    .io_b_6(dot_14_io_b_6),
    .io_b_7(dot_14_io_b_7),
    .io_b_8(dot_14_io_b_8),
    .io_b_9(dot_14_io_b_9),
    .io_b_10(dot_14_io_b_10),
    .io_b_11(dot_14_io_b_11),
    .io_b_12(dot_14_io_b_12),
    .io_b_13(dot_14_io_b_13),
    .io_b_14(dot_14_io_b_14),
    .io_b_15(dot_14_io_b_15),
    .io_y(dot_14_io_y)
  );
  DotProduct dot_15 ( // @[TensorGemm.scala 153:11:@18719.4]
    .clock(dot_15_clock),
    .io_a_0(dot_15_io_a_0),
    .io_a_1(dot_15_io_a_1),
    .io_a_2(dot_15_io_a_2),
    .io_a_3(dot_15_io_a_3),
    .io_a_4(dot_15_io_a_4),
    .io_a_5(dot_15_io_a_5),
    .io_a_6(dot_15_io_a_6),
    .io_a_7(dot_15_io_a_7),
    .io_a_8(dot_15_io_a_8),
    .io_a_9(dot_15_io_a_9),
    .io_a_10(dot_15_io_a_10),
    .io_a_11(dot_15_io_a_11),
    .io_a_12(dot_15_io_a_12),
    .io_a_13(dot_15_io_a_13),
    .io_a_14(dot_15_io_a_14),
    .io_a_15(dot_15_io_a_15),
    .io_b_0(dot_15_io_b_0),
    .io_b_1(dot_15_io_b_1),
    .io_b_2(dot_15_io_b_2),
    .io_b_3(dot_15_io_b_3),
    .io_b_4(dot_15_io_b_4),
    .io_b_5(dot_15_io_b_5),
    .io_b_6(dot_15_io_b_6),
    .io_b_7(dot_15_io_b_7),
    .io_b_8(dot_15_io_b_8),
    .io_b_9(dot_15_io_b_9),
    .io_b_10(dot_15_io_b_10),
    .io_b_11(dot_15_io_b_11),
    .io_b_12(dot_15_io_b_12),
    .io_b_13(dot_15_io_b_13),
    .io_b_14(dot_15_io_b_14),
    .io_b_15(dot_15_io_b_15),
    .io_y(dot_15_io_y)
  );
  Pipe acc_0 ( // @[TensorGemm.scala 156:34:@18722.4]
    .clock(acc_0_clock),
    .reset(acc_0_reset),
    .io_enq_valid(acc_0_io_enq_valid),
    .io_enq_bits(acc_0_io_enq_bits),
    .io_deq_valid(acc_0_io_deq_valid),
    .io_deq_bits(acc_0_io_deq_bits)
  );
  Pipe acc_1 ( // @[TensorGemm.scala 156:34:@18725.4]
    .clock(acc_1_clock),
    .reset(acc_1_reset),
    .io_enq_valid(acc_1_io_enq_valid),
    .io_enq_bits(acc_1_io_enq_bits),
    .io_deq_valid(acc_1_io_deq_valid),
    .io_deq_bits(acc_1_io_deq_bits)
  );
  Pipe acc_2 ( // @[TensorGemm.scala 156:34:@18728.4]
    .clock(acc_2_clock),
    .reset(acc_2_reset),
    .io_enq_valid(acc_2_io_enq_valid),
    .io_enq_bits(acc_2_io_enq_bits),
    .io_deq_valid(acc_2_io_deq_valid),
    .io_deq_bits(acc_2_io_deq_bits)
  );
  Pipe acc_3 ( // @[TensorGemm.scala 156:34:@18731.4]
    .clock(acc_3_clock),
    .reset(acc_3_reset),
    .io_enq_valid(acc_3_io_enq_valid),
    .io_enq_bits(acc_3_io_enq_bits),
    .io_deq_valid(acc_3_io_deq_valid),
    .io_deq_bits(acc_3_io_deq_bits)
  );
  Pipe acc_4 ( // @[TensorGemm.scala 156:34:@18734.4]
    .clock(acc_4_clock),
    .reset(acc_4_reset),
    .io_enq_valid(acc_4_io_enq_valid),
    .io_enq_bits(acc_4_io_enq_bits),
    .io_deq_valid(acc_4_io_deq_valid),
    .io_deq_bits(acc_4_io_deq_bits)
  );
  Pipe acc_5 ( // @[TensorGemm.scala 156:34:@18737.4]
    .clock(acc_5_clock),
    .reset(acc_5_reset),
    .io_enq_valid(acc_5_io_enq_valid),
    .io_enq_bits(acc_5_io_enq_bits),
    .io_deq_valid(acc_5_io_deq_valid),
    .io_deq_bits(acc_5_io_deq_bits)
  );
  Pipe acc_6 ( // @[TensorGemm.scala 156:34:@18740.4]
    .clock(acc_6_clock),
    .reset(acc_6_reset),
    .io_enq_valid(acc_6_io_enq_valid),
    .io_enq_bits(acc_6_io_enq_bits),
    .io_deq_valid(acc_6_io_deq_valid),
    .io_deq_bits(acc_6_io_deq_bits)
  );
  Pipe acc_7 ( // @[TensorGemm.scala 156:34:@18743.4]
    .clock(acc_7_clock),
    .reset(acc_7_reset),
    .io_enq_valid(acc_7_io_enq_valid),
    .io_enq_bits(acc_7_io_enq_bits),
    .io_deq_valid(acc_7_io_deq_valid),
    .io_deq_bits(acc_7_io_deq_bits)
  );
  Pipe acc_8 ( // @[TensorGemm.scala 156:34:@18746.4]
    .clock(acc_8_clock),
    .reset(acc_8_reset),
    .io_enq_valid(acc_8_io_enq_valid),
    .io_enq_bits(acc_8_io_enq_bits),
    .io_deq_valid(acc_8_io_deq_valid),
    .io_deq_bits(acc_8_io_deq_bits)
  );
  Pipe acc_9 ( // @[TensorGemm.scala 156:34:@18749.4]
    .clock(acc_9_clock),
    .reset(acc_9_reset),
    .io_enq_valid(acc_9_io_enq_valid),
    .io_enq_bits(acc_9_io_enq_bits),
    .io_deq_valid(acc_9_io_deq_valid),
    .io_deq_bits(acc_9_io_deq_bits)
  );
  Pipe acc_10 ( // @[TensorGemm.scala 156:34:@18752.4]
    .clock(acc_10_clock),
    .reset(acc_10_reset),
    .io_enq_valid(acc_10_io_enq_valid),
    .io_enq_bits(acc_10_io_enq_bits),
    .io_deq_valid(acc_10_io_deq_valid),
    .io_deq_bits(acc_10_io_deq_bits)
  );
  Pipe acc_11 ( // @[TensorGemm.scala 156:34:@18755.4]
    .clock(acc_11_clock),
    .reset(acc_11_reset),
    .io_enq_valid(acc_11_io_enq_valid),
    .io_enq_bits(acc_11_io_enq_bits),
    .io_deq_valid(acc_11_io_deq_valid),
    .io_deq_bits(acc_11_io_deq_bits)
  );
  Pipe acc_12 ( // @[TensorGemm.scala 156:34:@18758.4]
    .clock(acc_12_clock),
    .reset(acc_12_reset),
    .io_enq_valid(acc_12_io_enq_valid),
    .io_enq_bits(acc_12_io_enq_bits),
    .io_deq_valid(acc_12_io_deq_valid),
    .io_deq_bits(acc_12_io_deq_bits)
  );
  Pipe acc_13 ( // @[TensorGemm.scala 156:34:@18761.4]
    .clock(acc_13_clock),
    .reset(acc_13_reset),
    .io_enq_valid(acc_13_io_enq_valid),
    .io_enq_bits(acc_13_io_enq_bits),
    .io_deq_valid(acc_13_io_deq_valid),
    .io_deq_bits(acc_13_io_deq_bits)
  );
  Pipe acc_14 ( // @[TensorGemm.scala 156:34:@18764.4]
    .clock(acc_14_clock),
    .reset(acc_14_reset),
    .io_enq_valid(acc_14_io_enq_valid),
    .io_enq_bits(acc_14_io_enq_bits),
    .io_deq_valid(acc_14_io_deq_valid),
    .io_deq_bits(acc_14_io_deq_bits)
  );
  Pipe acc_15 ( // @[TensorGemm.scala 156:34:@18767.4]
    .clock(acc_15_clock),
    .reset(acc_15_reset),
    .io_enq_valid(acc_15_io_enq_valid),
    .io_enq_bits(acc_15_io_enq_bits),
    .io_deq_valid(acc_15_io_deq_valid),
    .io_deq_bits(acc_15_io_deq_bits)
  );
  assign _T_6016 = io_inp_data_valid & io_wgt_data_valid; // @[TensorGemm.scala 161:46:@18787.4]
  assign _T_6017 = _T_6016 & io_acc_i_data_valid; // @[TensorGemm.scala 161:66:@18788.4]
  assign _T_6018 = ~ io_reset; // @[TensorGemm.scala 161:90:@18789.4]
  assign _T_6052 = $signed(acc_0_io_deq_bits); // @[TensorGemm.scala 167:34:@18857.4]
  assign _GEN_0 = {{11{dot_0_io_y[20]}},dot_0_io_y}; // @[TensorGemm.scala 167:41:@18858.4]
  assign _T_6053 = $signed(_T_6052) + $signed(_GEN_0); // @[TensorGemm.scala 167:41:@18858.4]
  assign _T_6054 = $signed(_T_6052) + $signed(_GEN_0); // @[TensorGemm.scala 167:41:@18859.4]
  assign add_0 = $signed(_T_6054); // @[TensorGemm.scala 167:41:@18860.4]
  assign _T_6057 = $unsigned(add_0); // @[TensorGemm.scala 168:59:@18862.4]
  assign _T_6096 = $signed(acc_1_io_deq_bits); // @[TensorGemm.scala 167:34:@18938.4]
  assign _GEN_1 = {{11{dot_1_io_y[20]}},dot_1_io_y}; // @[TensorGemm.scala 167:41:@18939.4]
  assign _T_6097 = $signed(_T_6096) + $signed(_GEN_1); // @[TensorGemm.scala 167:41:@18939.4]
  assign _T_6098 = $signed(_T_6096) + $signed(_GEN_1); // @[TensorGemm.scala 167:41:@18940.4]
  assign add_1 = $signed(_T_6098); // @[TensorGemm.scala 167:41:@18941.4]
  assign _T_6101 = $unsigned(add_1); // @[TensorGemm.scala 168:59:@18943.4]
  assign _T_6140 = $signed(acc_2_io_deq_bits); // @[TensorGemm.scala 167:34:@19019.4]
  assign _GEN_2 = {{11{dot_2_io_y[20]}},dot_2_io_y}; // @[TensorGemm.scala 167:41:@19020.4]
  assign _T_6141 = $signed(_T_6140) + $signed(_GEN_2); // @[TensorGemm.scala 167:41:@19020.4]
  assign _T_6142 = $signed(_T_6140) + $signed(_GEN_2); // @[TensorGemm.scala 167:41:@19021.4]
  assign add_2 = $signed(_T_6142); // @[TensorGemm.scala 167:41:@19022.4]
  assign _T_6145 = $unsigned(add_2); // @[TensorGemm.scala 168:59:@19024.4]
  assign _T_6184 = $signed(acc_3_io_deq_bits); // @[TensorGemm.scala 167:34:@19100.4]
  assign _GEN_3 = {{11{dot_3_io_y[20]}},dot_3_io_y}; // @[TensorGemm.scala 167:41:@19101.4]
  assign _T_6185 = $signed(_T_6184) + $signed(_GEN_3); // @[TensorGemm.scala 167:41:@19101.4]
  assign _T_6186 = $signed(_T_6184) + $signed(_GEN_3); // @[TensorGemm.scala 167:41:@19102.4]
  assign add_3 = $signed(_T_6186); // @[TensorGemm.scala 167:41:@19103.4]
  assign _T_6189 = $unsigned(add_3); // @[TensorGemm.scala 168:59:@19105.4]
  assign _T_6228 = $signed(acc_4_io_deq_bits); // @[TensorGemm.scala 167:34:@19181.4]
  assign _GEN_4 = {{11{dot_4_io_y[20]}},dot_4_io_y}; // @[TensorGemm.scala 167:41:@19182.4]
  assign _T_6229 = $signed(_T_6228) + $signed(_GEN_4); // @[TensorGemm.scala 167:41:@19182.4]
  assign _T_6230 = $signed(_T_6228) + $signed(_GEN_4); // @[TensorGemm.scala 167:41:@19183.4]
  assign add_4 = $signed(_T_6230); // @[TensorGemm.scala 167:41:@19184.4]
  assign _T_6233 = $unsigned(add_4); // @[TensorGemm.scala 168:59:@19186.4]
  assign _T_6272 = $signed(acc_5_io_deq_bits); // @[TensorGemm.scala 167:34:@19262.4]
  assign _GEN_5 = {{11{dot_5_io_y[20]}},dot_5_io_y}; // @[TensorGemm.scala 167:41:@19263.4]
  assign _T_6273 = $signed(_T_6272) + $signed(_GEN_5); // @[TensorGemm.scala 167:41:@19263.4]
  assign _T_6274 = $signed(_T_6272) + $signed(_GEN_5); // @[TensorGemm.scala 167:41:@19264.4]
  assign add_5 = $signed(_T_6274); // @[TensorGemm.scala 167:41:@19265.4]
  assign _T_6277 = $unsigned(add_5); // @[TensorGemm.scala 168:59:@19267.4]
  assign _T_6316 = $signed(acc_6_io_deq_bits); // @[TensorGemm.scala 167:34:@19343.4]
  assign _GEN_6 = {{11{dot_6_io_y[20]}},dot_6_io_y}; // @[TensorGemm.scala 167:41:@19344.4]
  assign _T_6317 = $signed(_T_6316) + $signed(_GEN_6); // @[TensorGemm.scala 167:41:@19344.4]
  assign _T_6318 = $signed(_T_6316) + $signed(_GEN_6); // @[TensorGemm.scala 167:41:@19345.4]
  assign add_6 = $signed(_T_6318); // @[TensorGemm.scala 167:41:@19346.4]
  assign _T_6321 = $unsigned(add_6); // @[TensorGemm.scala 168:59:@19348.4]
  assign _T_6360 = $signed(acc_7_io_deq_bits); // @[TensorGemm.scala 167:34:@19424.4]
  assign _GEN_7 = {{11{dot_7_io_y[20]}},dot_7_io_y}; // @[TensorGemm.scala 167:41:@19425.4]
  assign _T_6361 = $signed(_T_6360) + $signed(_GEN_7); // @[TensorGemm.scala 167:41:@19425.4]
  assign _T_6362 = $signed(_T_6360) + $signed(_GEN_7); // @[TensorGemm.scala 167:41:@19426.4]
  assign add_7 = $signed(_T_6362); // @[TensorGemm.scala 167:41:@19427.4]
  assign _T_6365 = $unsigned(add_7); // @[TensorGemm.scala 168:59:@19429.4]
  assign _T_6404 = $signed(acc_8_io_deq_bits); // @[TensorGemm.scala 167:34:@19505.4]
  assign _GEN_8 = {{11{dot_8_io_y[20]}},dot_8_io_y}; // @[TensorGemm.scala 167:41:@19506.4]
  assign _T_6405 = $signed(_T_6404) + $signed(_GEN_8); // @[TensorGemm.scala 167:41:@19506.4]
  assign _T_6406 = $signed(_T_6404) + $signed(_GEN_8); // @[TensorGemm.scala 167:41:@19507.4]
  assign add_8 = $signed(_T_6406); // @[TensorGemm.scala 167:41:@19508.4]
  assign _T_6409 = $unsigned(add_8); // @[TensorGemm.scala 168:59:@19510.4]
  assign _T_6448 = $signed(acc_9_io_deq_bits); // @[TensorGemm.scala 167:34:@19586.4]
  assign _GEN_9 = {{11{dot_9_io_y[20]}},dot_9_io_y}; // @[TensorGemm.scala 167:41:@19587.4]
  assign _T_6449 = $signed(_T_6448) + $signed(_GEN_9); // @[TensorGemm.scala 167:41:@19587.4]
  assign _T_6450 = $signed(_T_6448) + $signed(_GEN_9); // @[TensorGemm.scala 167:41:@19588.4]
  assign add_9 = $signed(_T_6450); // @[TensorGemm.scala 167:41:@19589.4]
  assign _T_6453 = $unsigned(add_9); // @[TensorGemm.scala 168:59:@19591.4]
  assign _T_6492 = $signed(acc_10_io_deq_bits); // @[TensorGemm.scala 167:34:@19667.4]
  assign _GEN_10 = {{11{dot_10_io_y[20]}},dot_10_io_y}; // @[TensorGemm.scala 167:41:@19668.4]
  assign _T_6493 = $signed(_T_6492) + $signed(_GEN_10); // @[TensorGemm.scala 167:41:@19668.4]
  assign _T_6494 = $signed(_T_6492) + $signed(_GEN_10); // @[TensorGemm.scala 167:41:@19669.4]
  assign add_10 = $signed(_T_6494); // @[TensorGemm.scala 167:41:@19670.4]
  assign _T_6497 = $unsigned(add_10); // @[TensorGemm.scala 168:59:@19672.4]
  assign _T_6536 = $signed(acc_11_io_deq_bits); // @[TensorGemm.scala 167:34:@19748.4]
  assign _GEN_11 = {{11{dot_11_io_y[20]}},dot_11_io_y}; // @[TensorGemm.scala 167:41:@19749.4]
  assign _T_6537 = $signed(_T_6536) + $signed(_GEN_11); // @[TensorGemm.scala 167:41:@19749.4]
  assign _T_6538 = $signed(_T_6536) + $signed(_GEN_11); // @[TensorGemm.scala 167:41:@19750.4]
  assign add_11 = $signed(_T_6538); // @[TensorGemm.scala 167:41:@19751.4]
  assign _T_6541 = $unsigned(add_11); // @[TensorGemm.scala 168:59:@19753.4]
  assign _T_6580 = $signed(acc_12_io_deq_bits); // @[TensorGemm.scala 167:34:@19829.4]
  assign _GEN_12 = {{11{dot_12_io_y[20]}},dot_12_io_y}; // @[TensorGemm.scala 167:41:@19830.4]
  assign _T_6581 = $signed(_T_6580) + $signed(_GEN_12); // @[TensorGemm.scala 167:41:@19830.4]
  assign _T_6582 = $signed(_T_6580) + $signed(_GEN_12); // @[TensorGemm.scala 167:41:@19831.4]
  assign add_12 = $signed(_T_6582); // @[TensorGemm.scala 167:41:@19832.4]
  assign _T_6585 = $unsigned(add_12); // @[TensorGemm.scala 168:59:@19834.4]
  assign _T_6624 = $signed(acc_13_io_deq_bits); // @[TensorGemm.scala 167:34:@19910.4]
  assign _GEN_13 = {{11{dot_13_io_y[20]}},dot_13_io_y}; // @[TensorGemm.scala 167:41:@19911.4]
  assign _T_6625 = $signed(_T_6624) + $signed(_GEN_13); // @[TensorGemm.scala 167:41:@19911.4]
  assign _T_6626 = $signed(_T_6624) + $signed(_GEN_13); // @[TensorGemm.scala 167:41:@19912.4]
  assign add_13 = $signed(_T_6626); // @[TensorGemm.scala 167:41:@19913.4]
  assign _T_6629 = $unsigned(add_13); // @[TensorGemm.scala 168:59:@19915.4]
  assign _T_6668 = $signed(acc_14_io_deq_bits); // @[TensorGemm.scala 167:34:@19991.4]
  assign _GEN_14 = {{11{dot_14_io_y[20]}},dot_14_io_y}; // @[TensorGemm.scala 167:41:@19992.4]
  assign _T_6669 = $signed(_T_6668) + $signed(_GEN_14); // @[TensorGemm.scala 167:41:@19992.4]
  assign _T_6670 = $signed(_T_6668) + $signed(_GEN_14); // @[TensorGemm.scala 167:41:@19993.4]
  assign add_14 = $signed(_T_6670); // @[TensorGemm.scala 167:41:@19994.4]
  assign _T_6673 = $unsigned(add_14); // @[TensorGemm.scala 168:59:@19996.4]
  assign _T_6712 = $signed(acc_15_io_deq_bits); // @[TensorGemm.scala 167:34:@20072.4]
  assign _GEN_15 = {{11{dot_15_io_y[20]}},dot_15_io_y}; // @[TensorGemm.scala 167:41:@20073.4]
  assign _T_6713 = $signed(_T_6712) + $signed(_GEN_15); // @[TensorGemm.scala 167:41:@20073.4]
  assign _T_6714 = $signed(_T_6712) + $signed(_GEN_15); // @[TensorGemm.scala 167:41:@20074.4]
  assign add_15 = $signed(_T_6714); // @[TensorGemm.scala 167:41:@20075.4]
  assign _T_6717 = $unsigned(add_15); // @[TensorGemm.scala 168:59:@20077.4]
  assign vld_1 = acc_1_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@18948.4]
  assign vld_0 = acc_0_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@18867.4]
  assign vld_3 = acc_3_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19110.4]
  assign vld_2 = acc_2_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19029.4]
  assign vld_5 = acc_5_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19272.4]
  assign vld_4 = acc_4_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19191.4]
  assign vld_7 = acc_7_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19434.4]
  assign vld_6 = acc_6_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19353.4]
  assign _T_6726 = {vld_7,vld_6,vld_5,vld_4,vld_3,vld_2,vld_1,vld_0}; // @[TensorGemm.scala 172:30:@20089.4]
  assign vld_9 = acc_9_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19596.4]
  assign vld_8 = acc_8_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19515.4]
  assign vld_11 = acc_11_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19758.4]
  assign vld_10 = acc_10_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19677.4]
  assign vld_13 = acc_13_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19920.4]
  assign vld_12 = acc_12_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@19839.4]
  assign vld_15 = acc_15_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@20082.4]
  assign vld_14 = acc_14_io_deq_valid; // @[TensorGemm.scala 158:17:@18786.4 TensorGemm.scala 170:12:@20001.4]
  assign _T_6734 = {vld_15,vld_14,vld_13,vld_12,vld_11,vld_10,vld_9,vld_8,_T_6726}; // @[TensorGemm.scala 172:30:@20097.4]
  assign _T_6735 = ~ _T_6734; // @[TensorGemm.scala 172:37:@20098.4]
  assign _T_6737 = _T_6735 == 16'h0; // @[TensorGemm.scala 172:37:@20099.4]
  assign io_acc_o_data_valid = _T_6737 | io_reset; // @[TensorGemm.scala 172:23:@20101.4]
  assign io_acc_o_data_bits_0_0 = io_reset ? 32'h0 : _T_6057; // @[TensorGemm.scala 168:30:@18864.4]
  assign io_acc_o_data_bits_0_1 = io_reset ? 32'h0 : _T_6101; // @[TensorGemm.scala 168:30:@18945.4]
  assign io_acc_o_data_bits_0_2 = io_reset ? 32'h0 : _T_6145; // @[TensorGemm.scala 168:30:@19026.4]
  assign io_acc_o_data_bits_0_3 = io_reset ? 32'h0 : _T_6189; // @[TensorGemm.scala 168:30:@19107.4]
  assign io_acc_o_data_bits_0_4 = io_reset ? 32'h0 : _T_6233; // @[TensorGemm.scala 168:30:@19188.4]
  assign io_acc_o_data_bits_0_5 = io_reset ? 32'h0 : _T_6277; // @[TensorGemm.scala 168:30:@19269.4]
  assign io_acc_o_data_bits_0_6 = io_reset ? 32'h0 : _T_6321; // @[TensorGemm.scala 168:30:@19350.4]
  assign io_acc_o_data_bits_0_7 = io_reset ? 32'h0 : _T_6365; // @[TensorGemm.scala 168:30:@19431.4]
  assign io_acc_o_data_bits_0_8 = io_reset ? 32'h0 : _T_6409; // @[TensorGemm.scala 168:30:@19512.4]
  assign io_acc_o_data_bits_0_9 = io_reset ? 32'h0 : _T_6453; // @[TensorGemm.scala 168:30:@19593.4]
  assign io_acc_o_data_bits_0_10 = io_reset ? 32'h0 : _T_6497; // @[TensorGemm.scala 168:30:@19674.4]
  assign io_acc_o_data_bits_0_11 = io_reset ? 32'h0 : _T_6541; // @[TensorGemm.scala 168:30:@19755.4]
  assign io_acc_o_data_bits_0_12 = io_reset ? 32'h0 : _T_6585; // @[TensorGemm.scala 168:30:@19836.4]
  assign io_acc_o_data_bits_0_13 = io_reset ? 32'h0 : _T_6629; // @[TensorGemm.scala 168:30:@19917.4]
  assign io_acc_o_data_bits_0_14 = io_reset ? 32'h0 : _T_6673; // @[TensorGemm.scala 168:30:@19998.4]
  assign io_acc_o_data_bits_0_15 = io_reset ? 32'h0 : _T_6717; // @[TensorGemm.scala 168:30:@20079.4]
  assign io_out_data_valid = _T_6735 == 16'h0; // @[TensorGemm.scala 173:21:@20119.4]
  assign io_out_data_bits_0_0 = _T_6057[7:0]; // @[TensorGemm.scala 169:28:@18866.4]
  assign io_out_data_bits_0_1 = _T_6101[7:0]; // @[TensorGemm.scala 169:28:@18947.4]
  assign io_out_data_bits_0_2 = _T_6145[7:0]; // @[TensorGemm.scala 169:28:@19028.4]
  assign io_out_data_bits_0_3 = _T_6189[7:0]; // @[TensorGemm.scala 169:28:@19109.4]
  assign io_out_data_bits_0_4 = _T_6233[7:0]; // @[TensorGemm.scala 169:28:@19190.4]
  assign io_out_data_bits_0_5 = _T_6277[7:0]; // @[TensorGemm.scala 169:28:@19271.4]
  assign io_out_data_bits_0_6 = _T_6321[7:0]; // @[TensorGemm.scala 169:28:@19352.4]
  assign io_out_data_bits_0_7 = _T_6365[7:0]; // @[TensorGemm.scala 169:28:@19433.4]
  assign io_out_data_bits_0_8 = _T_6409[7:0]; // @[TensorGemm.scala 169:28:@19514.4]
  assign io_out_data_bits_0_9 = _T_6453[7:0]; // @[TensorGemm.scala 169:28:@19595.4]
  assign io_out_data_bits_0_10 = _T_6497[7:0]; // @[TensorGemm.scala 169:28:@19676.4]
  assign io_out_data_bits_0_11 = _T_6541[7:0]; // @[TensorGemm.scala 169:28:@19757.4]
  assign io_out_data_bits_0_12 = _T_6585[7:0]; // @[TensorGemm.scala 169:28:@19838.4]
  assign io_out_data_bits_0_13 = _T_6629[7:0]; // @[TensorGemm.scala 169:28:@19919.4]
  assign io_out_data_bits_0_14 = _T_6673[7:0]; // @[TensorGemm.scala 169:28:@20000.4]
  assign io_out_data_bits_0_15 = _T_6717[7:0]; // @[TensorGemm.scala 169:28:@20081.4]
  assign dot_0_clock = clock; // @[:@18675.4]
  assign dot_0_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@18794.4]
  assign dot_0_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@18798.4]
  assign dot_0_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@18802.4]
  assign dot_0_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@18806.4]
  assign dot_0_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@18810.4]
  assign dot_0_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@18814.4]
  assign dot_0_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@18818.4]
  assign dot_0_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@18822.4]
  assign dot_0_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@18826.4]
  assign dot_0_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@18830.4]
  assign dot_0_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@18834.4]
  assign dot_0_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@18838.4]
  assign dot_0_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@18842.4]
  assign dot_0_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@18846.4]
  assign dot_0_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@18850.4]
  assign dot_0_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@18854.4]
  assign dot_0_io_b_0 = $signed(io_wgt_data_bits_0_0); // @[TensorGemm.scala 165:22:@18796.4]
  assign dot_0_io_b_1 = $signed(io_wgt_data_bits_0_1); // @[TensorGemm.scala 165:22:@18800.4]
  assign dot_0_io_b_2 = $signed(io_wgt_data_bits_0_2); // @[TensorGemm.scala 165:22:@18804.4]
  assign dot_0_io_b_3 = $signed(io_wgt_data_bits_0_3); // @[TensorGemm.scala 165:22:@18808.4]
  assign dot_0_io_b_4 = $signed(io_wgt_data_bits_0_4); // @[TensorGemm.scala 165:22:@18812.4]
  assign dot_0_io_b_5 = $signed(io_wgt_data_bits_0_5); // @[TensorGemm.scala 165:22:@18816.4]
  assign dot_0_io_b_6 = $signed(io_wgt_data_bits_0_6); // @[TensorGemm.scala 165:22:@18820.4]
  assign dot_0_io_b_7 = $signed(io_wgt_data_bits_0_7); // @[TensorGemm.scala 165:22:@18824.4]
  assign dot_0_io_b_8 = $signed(io_wgt_data_bits_0_8); // @[TensorGemm.scala 165:22:@18828.4]
  assign dot_0_io_b_9 = $signed(io_wgt_data_bits_0_9); // @[TensorGemm.scala 165:22:@18832.4]
  assign dot_0_io_b_10 = $signed(io_wgt_data_bits_0_10); // @[TensorGemm.scala 165:22:@18836.4]
  assign dot_0_io_b_11 = $signed(io_wgt_data_bits_0_11); // @[TensorGemm.scala 165:22:@18840.4]
  assign dot_0_io_b_12 = $signed(io_wgt_data_bits_0_12); // @[TensorGemm.scala 165:22:@18844.4]
  assign dot_0_io_b_13 = $signed(io_wgt_data_bits_0_13); // @[TensorGemm.scala 165:22:@18848.4]
  assign dot_0_io_b_14 = $signed(io_wgt_data_bits_0_14); // @[TensorGemm.scala 165:22:@18852.4]
  assign dot_0_io_b_15 = $signed(io_wgt_data_bits_0_15); // @[TensorGemm.scala 165:22:@18856.4]
  assign dot_1_clock = clock; // @[:@18678.4]
  assign dot_1_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@18875.4]
  assign dot_1_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@18879.4]
  assign dot_1_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@18883.4]
  assign dot_1_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@18887.4]
  assign dot_1_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@18891.4]
  assign dot_1_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@18895.4]
  assign dot_1_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@18899.4]
  assign dot_1_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@18903.4]
  assign dot_1_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@18907.4]
  assign dot_1_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@18911.4]
  assign dot_1_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@18915.4]
  assign dot_1_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@18919.4]
  assign dot_1_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@18923.4]
  assign dot_1_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@18927.4]
  assign dot_1_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@18931.4]
  assign dot_1_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@18935.4]
  assign dot_1_io_b_0 = $signed(io_wgt_data_bits_1_0); // @[TensorGemm.scala 165:22:@18877.4]
  assign dot_1_io_b_1 = $signed(io_wgt_data_bits_1_1); // @[TensorGemm.scala 165:22:@18881.4]
  assign dot_1_io_b_2 = $signed(io_wgt_data_bits_1_2); // @[TensorGemm.scala 165:22:@18885.4]
  assign dot_1_io_b_3 = $signed(io_wgt_data_bits_1_3); // @[TensorGemm.scala 165:22:@18889.4]
  assign dot_1_io_b_4 = $signed(io_wgt_data_bits_1_4); // @[TensorGemm.scala 165:22:@18893.4]
  assign dot_1_io_b_5 = $signed(io_wgt_data_bits_1_5); // @[TensorGemm.scala 165:22:@18897.4]
  assign dot_1_io_b_6 = $signed(io_wgt_data_bits_1_6); // @[TensorGemm.scala 165:22:@18901.4]
  assign dot_1_io_b_7 = $signed(io_wgt_data_bits_1_7); // @[TensorGemm.scala 165:22:@18905.4]
  assign dot_1_io_b_8 = $signed(io_wgt_data_bits_1_8); // @[TensorGemm.scala 165:22:@18909.4]
  assign dot_1_io_b_9 = $signed(io_wgt_data_bits_1_9); // @[TensorGemm.scala 165:22:@18913.4]
  assign dot_1_io_b_10 = $signed(io_wgt_data_bits_1_10); // @[TensorGemm.scala 165:22:@18917.4]
  assign dot_1_io_b_11 = $signed(io_wgt_data_bits_1_11); // @[TensorGemm.scala 165:22:@18921.4]
  assign dot_1_io_b_12 = $signed(io_wgt_data_bits_1_12); // @[TensorGemm.scala 165:22:@18925.4]
  assign dot_1_io_b_13 = $signed(io_wgt_data_bits_1_13); // @[TensorGemm.scala 165:22:@18929.4]
  assign dot_1_io_b_14 = $signed(io_wgt_data_bits_1_14); // @[TensorGemm.scala 165:22:@18933.4]
  assign dot_1_io_b_15 = $signed(io_wgt_data_bits_1_15); // @[TensorGemm.scala 165:22:@18937.4]
  assign dot_2_clock = clock; // @[:@18681.4]
  assign dot_2_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@18956.4]
  assign dot_2_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@18960.4]
  assign dot_2_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@18964.4]
  assign dot_2_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@18968.4]
  assign dot_2_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@18972.4]
  assign dot_2_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@18976.4]
  assign dot_2_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@18980.4]
  assign dot_2_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@18984.4]
  assign dot_2_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@18988.4]
  assign dot_2_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@18992.4]
  assign dot_2_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@18996.4]
  assign dot_2_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19000.4]
  assign dot_2_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19004.4]
  assign dot_2_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19008.4]
  assign dot_2_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19012.4]
  assign dot_2_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19016.4]
  assign dot_2_io_b_0 = $signed(io_wgt_data_bits_2_0); // @[TensorGemm.scala 165:22:@18958.4]
  assign dot_2_io_b_1 = $signed(io_wgt_data_bits_2_1); // @[TensorGemm.scala 165:22:@18962.4]
  assign dot_2_io_b_2 = $signed(io_wgt_data_bits_2_2); // @[TensorGemm.scala 165:22:@18966.4]
  assign dot_2_io_b_3 = $signed(io_wgt_data_bits_2_3); // @[TensorGemm.scala 165:22:@18970.4]
  assign dot_2_io_b_4 = $signed(io_wgt_data_bits_2_4); // @[TensorGemm.scala 165:22:@18974.4]
  assign dot_2_io_b_5 = $signed(io_wgt_data_bits_2_5); // @[TensorGemm.scala 165:22:@18978.4]
  assign dot_2_io_b_6 = $signed(io_wgt_data_bits_2_6); // @[TensorGemm.scala 165:22:@18982.4]
  assign dot_2_io_b_7 = $signed(io_wgt_data_bits_2_7); // @[TensorGemm.scala 165:22:@18986.4]
  assign dot_2_io_b_8 = $signed(io_wgt_data_bits_2_8); // @[TensorGemm.scala 165:22:@18990.4]
  assign dot_2_io_b_9 = $signed(io_wgt_data_bits_2_9); // @[TensorGemm.scala 165:22:@18994.4]
  assign dot_2_io_b_10 = $signed(io_wgt_data_bits_2_10); // @[TensorGemm.scala 165:22:@18998.4]
  assign dot_2_io_b_11 = $signed(io_wgt_data_bits_2_11); // @[TensorGemm.scala 165:22:@19002.4]
  assign dot_2_io_b_12 = $signed(io_wgt_data_bits_2_12); // @[TensorGemm.scala 165:22:@19006.4]
  assign dot_2_io_b_13 = $signed(io_wgt_data_bits_2_13); // @[TensorGemm.scala 165:22:@19010.4]
  assign dot_2_io_b_14 = $signed(io_wgt_data_bits_2_14); // @[TensorGemm.scala 165:22:@19014.4]
  assign dot_2_io_b_15 = $signed(io_wgt_data_bits_2_15); // @[TensorGemm.scala 165:22:@19018.4]
  assign dot_3_clock = clock; // @[:@18684.4]
  assign dot_3_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19037.4]
  assign dot_3_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19041.4]
  assign dot_3_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19045.4]
  assign dot_3_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19049.4]
  assign dot_3_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19053.4]
  assign dot_3_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19057.4]
  assign dot_3_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19061.4]
  assign dot_3_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19065.4]
  assign dot_3_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19069.4]
  assign dot_3_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19073.4]
  assign dot_3_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19077.4]
  assign dot_3_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19081.4]
  assign dot_3_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19085.4]
  assign dot_3_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19089.4]
  assign dot_3_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19093.4]
  assign dot_3_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19097.4]
  assign dot_3_io_b_0 = $signed(io_wgt_data_bits_3_0); // @[TensorGemm.scala 165:22:@19039.4]
  assign dot_3_io_b_1 = $signed(io_wgt_data_bits_3_1); // @[TensorGemm.scala 165:22:@19043.4]
  assign dot_3_io_b_2 = $signed(io_wgt_data_bits_3_2); // @[TensorGemm.scala 165:22:@19047.4]
  assign dot_3_io_b_3 = $signed(io_wgt_data_bits_3_3); // @[TensorGemm.scala 165:22:@19051.4]
  assign dot_3_io_b_4 = $signed(io_wgt_data_bits_3_4); // @[TensorGemm.scala 165:22:@19055.4]
  assign dot_3_io_b_5 = $signed(io_wgt_data_bits_3_5); // @[TensorGemm.scala 165:22:@19059.4]
  assign dot_3_io_b_6 = $signed(io_wgt_data_bits_3_6); // @[TensorGemm.scala 165:22:@19063.4]
  assign dot_3_io_b_7 = $signed(io_wgt_data_bits_3_7); // @[TensorGemm.scala 165:22:@19067.4]
  assign dot_3_io_b_8 = $signed(io_wgt_data_bits_3_8); // @[TensorGemm.scala 165:22:@19071.4]
  assign dot_3_io_b_9 = $signed(io_wgt_data_bits_3_9); // @[TensorGemm.scala 165:22:@19075.4]
  assign dot_3_io_b_10 = $signed(io_wgt_data_bits_3_10); // @[TensorGemm.scala 165:22:@19079.4]
  assign dot_3_io_b_11 = $signed(io_wgt_data_bits_3_11); // @[TensorGemm.scala 165:22:@19083.4]
  assign dot_3_io_b_12 = $signed(io_wgt_data_bits_3_12); // @[TensorGemm.scala 165:22:@19087.4]
  assign dot_3_io_b_13 = $signed(io_wgt_data_bits_3_13); // @[TensorGemm.scala 165:22:@19091.4]
  assign dot_3_io_b_14 = $signed(io_wgt_data_bits_3_14); // @[TensorGemm.scala 165:22:@19095.4]
  assign dot_3_io_b_15 = $signed(io_wgt_data_bits_3_15); // @[TensorGemm.scala 165:22:@19099.4]
  assign dot_4_clock = clock; // @[:@18687.4]
  assign dot_4_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19118.4]
  assign dot_4_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19122.4]
  assign dot_4_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19126.4]
  assign dot_4_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19130.4]
  assign dot_4_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19134.4]
  assign dot_4_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19138.4]
  assign dot_4_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19142.4]
  assign dot_4_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19146.4]
  assign dot_4_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19150.4]
  assign dot_4_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19154.4]
  assign dot_4_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19158.4]
  assign dot_4_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19162.4]
  assign dot_4_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19166.4]
  assign dot_4_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19170.4]
  assign dot_4_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19174.4]
  assign dot_4_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19178.4]
  assign dot_4_io_b_0 = $signed(io_wgt_data_bits_4_0); // @[TensorGemm.scala 165:22:@19120.4]
  assign dot_4_io_b_1 = $signed(io_wgt_data_bits_4_1); // @[TensorGemm.scala 165:22:@19124.4]
  assign dot_4_io_b_2 = $signed(io_wgt_data_bits_4_2); // @[TensorGemm.scala 165:22:@19128.4]
  assign dot_4_io_b_3 = $signed(io_wgt_data_bits_4_3); // @[TensorGemm.scala 165:22:@19132.4]
  assign dot_4_io_b_4 = $signed(io_wgt_data_bits_4_4); // @[TensorGemm.scala 165:22:@19136.4]
  assign dot_4_io_b_5 = $signed(io_wgt_data_bits_4_5); // @[TensorGemm.scala 165:22:@19140.4]
  assign dot_4_io_b_6 = $signed(io_wgt_data_bits_4_6); // @[TensorGemm.scala 165:22:@19144.4]
  assign dot_4_io_b_7 = $signed(io_wgt_data_bits_4_7); // @[TensorGemm.scala 165:22:@19148.4]
  assign dot_4_io_b_8 = $signed(io_wgt_data_bits_4_8); // @[TensorGemm.scala 165:22:@19152.4]
  assign dot_4_io_b_9 = $signed(io_wgt_data_bits_4_9); // @[TensorGemm.scala 165:22:@19156.4]
  assign dot_4_io_b_10 = $signed(io_wgt_data_bits_4_10); // @[TensorGemm.scala 165:22:@19160.4]
  assign dot_4_io_b_11 = $signed(io_wgt_data_bits_4_11); // @[TensorGemm.scala 165:22:@19164.4]
  assign dot_4_io_b_12 = $signed(io_wgt_data_bits_4_12); // @[TensorGemm.scala 165:22:@19168.4]
  assign dot_4_io_b_13 = $signed(io_wgt_data_bits_4_13); // @[TensorGemm.scala 165:22:@19172.4]
  assign dot_4_io_b_14 = $signed(io_wgt_data_bits_4_14); // @[TensorGemm.scala 165:22:@19176.4]
  assign dot_4_io_b_15 = $signed(io_wgt_data_bits_4_15); // @[TensorGemm.scala 165:22:@19180.4]
  assign dot_5_clock = clock; // @[:@18690.4]
  assign dot_5_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19199.4]
  assign dot_5_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19203.4]
  assign dot_5_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19207.4]
  assign dot_5_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19211.4]
  assign dot_5_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19215.4]
  assign dot_5_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19219.4]
  assign dot_5_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19223.4]
  assign dot_5_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19227.4]
  assign dot_5_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19231.4]
  assign dot_5_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19235.4]
  assign dot_5_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19239.4]
  assign dot_5_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19243.4]
  assign dot_5_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19247.4]
  assign dot_5_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19251.4]
  assign dot_5_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19255.4]
  assign dot_5_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19259.4]
  assign dot_5_io_b_0 = $signed(io_wgt_data_bits_5_0); // @[TensorGemm.scala 165:22:@19201.4]
  assign dot_5_io_b_1 = $signed(io_wgt_data_bits_5_1); // @[TensorGemm.scala 165:22:@19205.4]
  assign dot_5_io_b_2 = $signed(io_wgt_data_bits_5_2); // @[TensorGemm.scala 165:22:@19209.4]
  assign dot_5_io_b_3 = $signed(io_wgt_data_bits_5_3); // @[TensorGemm.scala 165:22:@19213.4]
  assign dot_5_io_b_4 = $signed(io_wgt_data_bits_5_4); // @[TensorGemm.scala 165:22:@19217.4]
  assign dot_5_io_b_5 = $signed(io_wgt_data_bits_5_5); // @[TensorGemm.scala 165:22:@19221.4]
  assign dot_5_io_b_6 = $signed(io_wgt_data_bits_5_6); // @[TensorGemm.scala 165:22:@19225.4]
  assign dot_5_io_b_7 = $signed(io_wgt_data_bits_5_7); // @[TensorGemm.scala 165:22:@19229.4]
  assign dot_5_io_b_8 = $signed(io_wgt_data_bits_5_8); // @[TensorGemm.scala 165:22:@19233.4]
  assign dot_5_io_b_9 = $signed(io_wgt_data_bits_5_9); // @[TensorGemm.scala 165:22:@19237.4]
  assign dot_5_io_b_10 = $signed(io_wgt_data_bits_5_10); // @[TensorGemm.scala 165:22:@19241.4]
  assign dot_5_io_b_11 = $signed(io_wgt_data_bits_5_11); // @[TensorGemm.scala 165:22:@19245.4]
  assign dot_5_io_b_12 = $signed(io_wgt_data_bits_5_12); // @[TensorGemm.scala 165:22:@19249.4]
  assign dot_5_io_b_13 = $signed(io_wgt_data_bits_5_13); // @[TensorGemm.scala 165:22:@19253.4]
  assign dot_5_io_b_14 = $signed(io_wgt_data_bits_5_14); // @[TensorGemm.scala 165:22:@19257.4]
  assign dot_5_io_b_15 = $signed(io_wgt_data_bits_5_15); // @[TensorGemm.scala 165:22:@19261.4]
  assign dot_6_clock = clock; // @[:@18693.4]
  assign dot_6_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19280.4]
  assign dot_6_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19284.4]
  assign dot_6_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19288.4]
  assign dot_6_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19292.4]
  assign dot_6_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19296.4]
  assign dot_6_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19300.4]
  assign dot_6_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19304.4]
  assign dot_6_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19308.4]
  assign dot_6_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19312.4]
  assign dot_6_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19316.4]
  assign dot_6_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19320.4]
  assign dot_6_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19324.4]
  assign dot_6_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19328.4]
  assign dot_6_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19332.4]
  assign dot_6_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19336.4]
  assign dot_6_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19340.4]
  assign dot_6_io_b_0 = $signed(io_wgt_data_bits_6_0); // @[TensorGemm.scala 165:22:@19282.4]
  assign dot_6_io_b_1 = $signed(io_wgt_data_bits_6_1); // @[TensorGemm.scala 165:22:@19286.4]
  assign dot_6_io_b_2 = $signed(io_wgt_data_bits_6_2); // @[TensorGemm.scala 165:22:@19290.4]
  assign dot_6_io_b_3 = $signed(io_wgt_data_bits_6_3); // @[TensorGemm.scala 165:22:@19294.4]
  assign dot_6_io_b_4 = $signed(io_wgt_data_bits_6_4); // @[TensorGemm.scala 165:22:@19298.4]
  assign dot_6_io_b_5 = $signed(io_wgt_data_bits_6_5); // @[TensorGemm.scala 165:22:@19302.4]
  assign dot_6_io_b_6 = $signed(io_wgt_data_bits_6_6); // @[TensorGemm.scala 165:22:@19306.4]
  assign dot_6_io_b_7 = $signed(io_wgt_data_bits_6_7); // @[TensorGemm.scala 165:22:@19310.4]
  assign dot_6_io_b_8 = $signed(io_wgt_data_bits_6_8); // @[TensorGemm.scala 165:22:@19314.4]
  assign dot_6_io_b_9 = $signed(io_wgt_data_bits_6_9); // @[TensorGemm.scala 165:22:@19318.4]
  assign dot_6_io_b_10 = $signed(io_wgt_data_bits_6_10); // @[TensorGemm.scala 165:22:@19322.4]
  assign dot_6_io_b_11 = $signed(io_wgt_data_bits_6_11); // @[TensorGemm.scala 165:22:@19326.4]
  assign dot_6_io_b_12 = $signed(io_wgt_data_bits_6_12); // @[TensorGemm.scala 165:22:@19330.4]
  assign dot_6_io_b_13 = $signed(io_wgt_data_bits_6_13); // @[TensorGemm.scala 165:22:@19334.4]
  assign dot_6_io_b_14 = $signed(io_wgt_data_bits_6_14); // @[TensorGemm.scala 165:22:@19338.4]
  assign dot_6_io_b_15 = $signed(io_wgt_data_bits_6_15); // @[TensorGemm.scala 165:22:@19342.4]
  assign dot_7_clock = clock; // @[:@18696.4]
  assign dot_7_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19361.4]
  assign dot_7_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19365.4]
  assign dot_7_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19369.4]
  assign dot_7_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19373.4]
  assign dot_7_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19377.4]
  assign dot_7_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19381.4]
  assign dot_7_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19385.4]
  assign dot_7_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19389.4]
  assign dot_7_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19393.4]
  assign dot_7_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19397.4]
  assign dot_7_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19401.4]
  assign dot_7_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19405.4]
  assign dot_7_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19409.4]
  assign dot_7_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19413.4]
  assign dot_7_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19417.4]
  assign dot_7_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19421.4]
  assign dot_7_io_b_0 = $signed(io_wgt_data_bits_7_0); // @[TensorGemm.scala 165:22:@19363.4]
  assign dot_7_io_b_1 = $signed(io_wgt_data_bits_7_1); // @[TensorGemm.scala 165:22:@19367.4]
  assign dot_7_io_b_2 = $signed(io_wgt_data_bits_7_2); // @[TensorGemm.scala 165:22:@19371.4]
  assign dot_7_io_b_3 = $signed(io_wgt_data_bits_7_3); // @[TensorGemm.scala 165:22:@19375.4]
  assign dot_7_io_b_4 = $signed(io_wgt_data_bits_7_4); // @[TensorGemm.scala 165:22:@19379.4]
  assign dot_7_io_b_5 = $signed(io_wgt_data_bits_7_5); // @[TensorGemm.scala 165:22:@19383.4]
  assign dot_7_io_b_6 = $signed(io_wgt_data_bits_7_6); // @[TensorGemm.scala 165:22:@19387.4]
  assign dot_7_io_b_7 = $signed(io_wgt_data_bits_7_7); // @[TensorGemm.scala 165:22:@19391.4]
  assign dot_7_io_b_8 = $signed(io_wgt_data_bits_7_8); // @[TensorGemm.scala 165:22:@19395.4]
  assign dot_7_io_b_9 = $signed(io_wgt_data_bits_7_9); // @[TensorGemm.scala 165:22:@19399.4]
  assign dot_7_io_b_10 = $signed(io_wgt_data_bits_7_10); // @[TensorGemm.scala 165:22:@19403.4]
  assign dot_7_io_b_11 = $signed(io_wgt_data_bits_7_11); // @[TensorGemm.scala 165:22:@19407.4]
  assign dot_7_io_b_12 = $signed(io_wgt_data_bits_7_12); // @[TensorGemm.scala 165:22:@19411.4]
  assign dot_7_io_b_13 = $signed(io_wgt_data_bits_7_13); // @[TensorGemm.scala 165:22:@19415.4]
  assign dot_7_io_b_14 = $signed(io_wgt_data_bits_7_14); // @[TensorGemm.scala 165:22:@19419.4]
  assign dot_7_io_b_15 = $signed(io_wgt_data_bits_7_15); // @[TensorGemm.scala 165:22:@19423.4]
  assign dot_8_clock = clock; // @[:@18699.4]
  assign dot_8_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19442.4]
  assign dot_8_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19446.4]
  assign dot_8_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19450.4]
  assign dot_8_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19454.4]
  assign dot_8_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19458.4]
  assign dot_8_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19462.4]
  assign dot_8_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19466.4]
  assign dot_8_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19470.4]
  assign dot_8_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19474.4]
  assign dot_8_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19478.4]
  assign dot_8_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19482.4]
  assign dot_8_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19486.4]
  assign dot_8_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19490.4]
  assign dot_8_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19494.4]
  assign dot_8_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19498.4]
  assign dot_8_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19502.4]
  assign dot_8_io_b_0 = $signed(io_wgt_data_bits_8_0); // @[TensorGemm.scala 165:22:@19444.4]
  assign dot_8_io_b_1 = $signed(io_wgt_data_bits_8_1); // @[TensorGemm.scala 165:22:@19448.4]
  assign dot_8_io_b_2 = $signed(io_wgt_data_bits_8_2); // @[TensorGemm.scala 165:22:@19452.4]
  assign dot_8_io_b_3 = $signed(io_wgt_data_bits_8_3); // @[TensorGemm.scala 165:22:@19456.4]
  assign dot_8_io_b_4 = $signed(io_wgt_data_bits_8_4); // @[TensorGemm.scala 165:22:@19460.4]
  assign dot_8_io_b_5 = $signed(io_wgt_data_bits_8_5); // @[TensorGemm.scala 165:22:@19464.4]
  assign dot_8_io_b_6 = $signed(io_wgt_data_bits_8_6); // @[TensorGemm.scala 165:22:@19468.4]
  assign dot_8_io_b_7 = $signed(io_wgt_data_bits_8_7); // @[TensorGemm.scala 165:22:@19472.4]
  assign dot_8_io_b_8 = $signed(io_wgt_data_bits_8_8); // @[TensorGemm.scala 165:22:@19476.4]
  assign dot_8_io_b_9 = $signed(io_wgt_data_bits_8_9); // @[TensorGemm.scala 165:22:@19480.4]
  assign dot_8_io_b_10 = $signed(io_wgt_data_bits_8_10); // @[TensorGemm.scala 165:22:@19484.4]
  assign dot_8_io_b_11 = $signed(io_wgt_data_bits_8_11); // @[TensorGemm.scala 165:22:@19488.4]
  assign dot_8_io_b_12 = $signed(io_wgt_data_bits_8_12); // @[TensorGemm.scala 165:22:@19492.4]
  assign dot_8_io_b_13 = $signed(io_wgt_data_bits_8_13); // @[TensorGemm.scala 165:22:@19496.4]
  assign dot_8_io_b_14 = $signed(io_wgt_data_bits_8_14); // @[TensorGemm.scala 165:22:@19500.4]
  assign dot_8_io_b_15 = $signed(io_wgt_data_bits_8_15); // @[TensorGemm.scala 165:22:@19504.4]
  assign dot_9_clock = clock; // @[:@18702.4]
  assign dot_9_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19523.4]
  assign dot_9_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19527.4]
  assign dot_9_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19531.4]
  assign dot_9_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19535.4]
  assign dot_9_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19539.4]
  assign dot_9_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19543.4]
  assign dot_9_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19547.4]
  assign dot_9_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19551.4]
  assign dot_9_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19555.4]
  assign dot_9_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19559.4]
  assign dot_9_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19563.4]
  assign dot_9_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19567.4]
  assign dot_9_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19571.4]
  assign dot_9_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19575.4]
  assign dot_9_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19579.4]
  assign dot_9_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19583.4]
  assign dot_9_io_b_0 = $signed(io_wgt_data_bits_9_0); // @[TensorGemm.scala 165:22:@19525.4]
  assign dot_9_io_b_1 = $signed(io_wgt_data_bits_9_1); // @[TensorGemm.scala 165:22:@19529.4]
  assign dot_9_io_b_2 = $signed(io_wgt_data_bits_9_2); // @[TensorGemm.scala 165:22:@19533.4]
  assign dot_9_io_b_3 = $signed(io_wgt_data_bits_9_3); // @[TensorGemm.scala 165:22:@19537.4]
  assign dot_9_io_b_4 = $signed(io_wgt_data_bits_9_4); // @[TensorGemm.scala 165:22:@19541.4]
  assign dot_9_io_b_5 = $signed(io_wgt_data_bits_9_5); // @[TensorGemm.scala 165:22:@19545.4]
  assign dot_9_io_b_6 = $signed(io_wgt_data_bits_9_6); // @[TensorGemm.scala 165:22:@19549.4]
  assign dot_9_io_b_7 = $signed(io_wgt_data_bits_9_7); // @[TensorGemm.scala 165:22:@19553.4]
  assign dot_9_io_b_8 = $signed(io_wgt_data_bits_9_8); // @[TensorGemm.scala 165:22:@19557.4]
  assign dot_9_io_b_9 = $signed(io_wgt_data_bits_9_9); // @[TensorGemm.scala 165:22:@19561.4]
  assign dot_9_io_b_10 = $signed(io_wgt_data_bits_9_10); // @[TensorGemm.scala 165:22:@19565.4]
  assign dot_9_io_b_11 = $signed(io_wgt_data_bits_9_11); // @[TensorGemm.scala 165:22:@19569.4]
  assign dot_9_io_b_12 = $signed(io_wgt_data_bits_9_12); // @[TensorGemm.scala 165:22:@19573.4]
  assign dot_9_io_b_13 = $signed(io_wgt_data_bits_9_13); // @[TensorGemm.scala 165:22:@19577.4]
  assign dot_9_io_b_14 = $signed(io_wgt_data_bits_9_14); // @[TensorGemm.scala 165:22:@19581.4]
  assign dot_9_io_b_15 = $signed(io_wgt_data_bits_9_15); // @[TensorGemm.scala 165:22:@19585.4]
  assign dot_10_clock = clock; // @[:@18705.4]
  assign dot_10_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19604.4]
  assign dot_10_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19608.4]
  assign dot_10_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19612.4]
  assign dot_10_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19616.4]
  assign dot_10_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19620.4]
  assign dot_10_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19624.4]
  assign dot_10_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19628.4]
  assign dot_10_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19632.4]
  assign dot_10_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19636.4]
  assign dot_10_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19640.4]
  assign dot_10_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19644.4]
  assign dot_10_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19648.4]
  assign dot_10_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19652.4]
  assign dot_10_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19656.4]
  assign dot_10_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19660.4]
  assign dot_10_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19664.4]
  assign dot_10_io_b_0 = $signed(io_wgt_data_bits_10_0); // @[TensorGemm.scala 165:22:@19606.4]
  assign dot_10_io_b_1 = $signed(io_wgt_data_bits_10_1); // @[TensorGemm.scala 165:22:@19610.4]
  assign dot_10_io_b_2 = $signed(io_wgt_data_bits_10_2); // @[TensorGemm.scala 165:22:@19614.4]
  assign dot_10_io_b_3 = $signed(io_wgt_data_bits_10_3); // @[TensorGemm.scala 165:22:@19618.4]
  assign dot_10_io_b_4 = $signed(io_wgt_data_bits_10_4); // @[TensorGemm.scala 165:22:@19622.4]
  assign dot_10_io_b_5 = $signed(io_wgt_data_bits_10_5); // @[TensorGemm.scala 165:22:@19626.4]
  assign dot_10_io_b_6 = $signed(io_wgt_data_bits_10_6); // @[TensorGemm.scala 165:22:@19630.4]
  assign dot_10_io_b_7 = $signed(io_wgt_data_bits_10_7); // @[TensorGemm.scala 165:22:@19634.4]
  assign dot_10_io_b_8 = $signed(io_wgt_data_bits_10_8); // @[TensorGemm.scala 165:22:@19638.4]
  assign dot_10_io_b_9 = $signed(io_wgt_data_bits_10_9); // @[TensorGemm.scala 165:22:@19642.4]
  assign dot_10_io_b_10 = $signed(io_wgt_data_bits_10_10); // @[TensorGemm.scala 165:22:@19646.4]
  assign dot_10_io_b_11 = $signed(io_wgt_data_bits_10_11); // @[TensorGemm.scala 165:22:@19650.4]
  assign dot_10_io_b_12 = $signed(io_wgt_data_bits_10_12); // @[TensorGemm.scala 165:22:@19654.4]
  assign dot_10_io_b_13 = $signed(io_wgt_data_bits_10_13); // @[TensorGemm.scala 165:22:@19658.4]
  assign dot_10_io_b_14 = $signed(io_wgt_data_bits_10_14); // @[TensorGemm.scala 165:22:@19662.4]
  assign dot_10_io_b_15 = $signed(io_wgt_data_bits_10_15); // @[TensorGemm.scala 165:22:@19666.4]
  assign dot_11_clock = clock; // @[:@18708.4]
  assign dot_11_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19685.4]
  assign dot_11_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19689.4]
  assign dot_11_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19693.4]
  assign dot_11_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19697.4]
  assign dot_11_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19701.4]
  assign dot_11_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19705.4]
  assign dot_11_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19709.4]
  assign dot_11_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19713.4]
  assign dot_11_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19717.4]
  assign dot_11_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19721.4]
  assign dot_11_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19725.4]
  assign dot_11_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19729.4]
  assign dot_11_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19733.4]
  assign dot_11_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19737.4]
  assign dot_11_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19741.4]
  assign dot_11_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19745.4]
  assign dot_11_io_b_0 = $signed(io_wgt_data_bits_11_0); // @[TensorGemm.scala 165:22:@19687.4]
  assign dot_11_io_b_1 = $signed(io_wgt_data_bits_11_1); // @[TensorGemm.scala 165:22:@19691.4]
  assign dot_11_io_b_2 = $signed(io_wgt_data_bits_11_2); // @[TensorGemm.scala 165:22:@19695.4]
  assign dot_11_io_b_3 = $signed(io_wgt_data_bits_11_3); // @[TensorGemm.scala 165:22:@19699.4]
  assign dot_11_io_b_4 = $signed(io_wgt_data_bits_11_4); // @[TensorGemm.scala 165:22:@19703.4]
  assign dot_11_io_b_5 = $signed(io_wgt_data_bits_11_5); // @[TensorGemm.scala 165:22:@19707.4]
  assign dot_11_io_b_6 = $signed(io_wgt_data_bits_11_6); // @[TensorGemm.scala 165:22:@19711.4]
  assign dot_11_io_b_7 = $signed(io_wgt_data_bits_11_7); // @[TensorGemm.scala 165:22:@19715.4]
  assign dot_11_io_b_8 = $signed(io_wgt_data_bits_11_8); // @[TensorGemm.scala 165:22:@19719.4]
  assign dot_11_io_b_9 = $signed(io_wgt_data_bits_11_9); // @[TensorGemm.scala 165:22:@19723.4]
  assign dot_11_io_b_10 = $signed(io_wgt_data_bits_11_10); // @[TensorGemm.scala 165:22:@19727.4]
  assign dot_11_io_b_11 = $signed(io_wgt_data_bits_11_11); // @[TensorGemm.scala 165:22:@19731.4]
  assign dot_11_io_b_12 = $signed(io_wgt_data_bits_11_12); // @[TensorGemm.scala 165:22:@19735.4]
  assign dot_11_io_b_13 = $signed(io_wgt_data_bits_11_13); // @[TensorGemm.scala 165:22:@19739.4]
  assign dot_11_io_b_14 = $signed(io_wgt_data_bits_11_14); // @[TensorGemm.scala 165:22:@19743.4]
  assign dot_11_io_b_15 = $signed(io_wgt_data_bits_11_15); // @[TensorGemm.scala 165:22:@19747.4]
  assign dot_12_clock = clock; // @[:@18711.4]
  assign dot_12_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19766.4]
  assign dot_12_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19770.4]
  assign dot_12_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19774.4]
  assign dot_12_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19778.4]
  assign dot_12_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19782.4]
  assign dot_12_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19786.4]
  assign dot_12_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19790.4]
  assign dot_12_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19794.4]
  assign dot_12_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19798.4]
  assign dot_12_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19802.4]
  assign dot_12_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19806.4]
  assign dot_12_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19810.4]
  assign dot_12_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19814.4]
  assign dot_12_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19818.4]
  assign dot_12_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19822.4]
  assign dot_12_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19826.4]
  assign dot_12_io_b_0 = $signed(io_wgt_data_bits_12_0); // @[TensorGemm.scala 165:22:@19768.4]
  assign dot_12_io_b_1 = $signed(io_wgt_data_bits_12_1); // @[TensorGemm.scala 165:22:@19772.4]
  assign dot_12_io_b_2 = $signed(io_wgt_data_bits_12_2); // @[TensorGemm.scala 165:22:@19776.4]
  assign dot_12_io_b_3 = $signed(io_wgt_data_bits_12_3); // @[TensorGemm.scala 165:22:@19780.4]
  assign dot_12_io_b_4 = $signed(io_wgt_data_bits_12_4); // @[TensorGemm.scala 165:22:@19784.4]
  assign dot_12_io_b_5 = $signed(io_wgt_data_bits_12_5); // @[TensorGemm.scala 165:22:@19788.4]
  assign dot_12_io_b_6 = $signed(io_wgt_data_bits_12_6); // @[TensorGemm.scala 165:22:@19792.4]
  assign dot_12_io_b_7 = $signed(io_wgt_data_bits_12_7); // @[TensorGemm.scala 165:22:@19796.4]
  assign dot_12_io_b_8 = $signed(io_wgt_data_bits_12_8); // @[TensorGemm.scala 165:22:@19800.4]
  assign dot_12_io_b_9 = $signed(io_wgt_data_bits_12_9); // @[TensorGemm.scala 165:22:@19804.4]
  assign dot_12_io_b_10 = $signed(io_wgt_data_bits_12_10); // @[TensorGemm.scala 165:22:@19808.4]
  assign dot_12_io_b_11 = $signed(io_wgt_data_bits_12_11); // @[TensorGemm.scala 165:22:@19812.4]
  assign dot_12_io_b_12 = $signed(io_wgt_data_bits_12_12); // @[TensorGemm.scala 165:22:@19816.4]
  assign dot_12_io_b_13 = $signed(io_wgt_data_bits_12_13); // @[TensorGemm.scala 165:22:@19820.4]
  assign dot_12_io_b_14 = $signed(io_wgt_data_bits_12_14); // @[TensorGemm.scala 165:22:@19824.4]
  assign dot_12_io_b_15 = $signed(io_wgt_data_bits_12_15); // @[TensorGemm.scala 165:22:@19828.4]
  assign dot_13_clock = clock; // @[:@18714.4]
  assign dot_13_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19847.4]
  assign dot_13_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19851.4]
  assign dot_13_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19855.4]
  assign dot_13_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19859.4]
  assign dot_13_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19863.4]
  assign dot_13_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19867.4]
  assign dot_13_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19871.4]
  assign dot_13_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19875.4]
  assign dot_13_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19879.4]
  assign dot_13_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19883.4]
  assign dot_13_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19887.4]
  assign dot_13_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19891.4]
  assign dot_13_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19895.4]
  assign dot_13_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19899.4]
  assign dot_13_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19903.4]
  assign dot_13_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19907.4]
  assign dot_13_io_b_0 = $signed(io_wgt_data_bits_13_0); // @[TensorGemm.scala 165:22:@19849.4]
  assign dot_13_io_b_1 = $signed(io_wgt_data_bits_13_1); // @[TensorGemm.scala 165:22:@19853.4]
  assign dot_13_io_b_2 = $signed(io_wgt_data_bits_13_2); // @[TensorGemm.scala 165:22:@19857.4]
  assign dot_13_io_b_3 = $signed(io_wgt_data_bits_13_3); // @[TensorGemm.scala 165:22:@19861.4]
  assign dot_13_io_b_4 = $signed(io_wgt_data_bits_13_4); // @[TensorGemm.scala 165:22:@19865.4]
  assign dot_13_io_b_5 = $signed(io_wgt_data_bits_13_5); // @[TensorGemm.scala 165:22:@19869.4]
  assign dot_13_io_b_6 = $signed(io_wgt_data_bits_13_6); // @[TensorGemm.scala 165:22:@19873.4]
  assign dot_13_io_b_7 = $signed(io_wgt_data_bits_13_7); // @[TensorGemm.scala 165:22:@19877.4]
  assign dot_13_io_b_8 = $signed(io_wgt_data_bits_13_8); // @[TensorGemm.scala 165:22:@19881.4]
  assign dot_13_io_b_9 = $signed(io_wgt_data_bits_13_9); // @[TensorGemm.scala 165:22:@19885.4]
  assign dot_13_io_b_10 = $signed(io_wgt_data_bits_13_10); // @[TensorGemm.scala 165:22:@19889.4]
  assign dot_13_io_b_11 = $signed(io_wgt_data_bits_13_11); // @[TensorGemm.scala 165:22:@19893.4]
  assign dot_13_io_b_12 = $signed(io_wgt_data_bits_13_12); // @[TensorGemm.scala 165:22:@19897.4]
  assign dot_13_io_b_13 = $signed(io_wgt_data_bits_13_13); // @[TensorGemm.scala 165:22:@19901.4]
  assign dot_13_io_b_14 = $signed(io_wgt_data_bits_13_14); // @[TensorGemm.scala 165:22:@19905.4]
  assign dot_13_io_b_15 = $signed(io_wgt_data_bits_13_15); // @[TensorGemm.scala 165:22:@19909.4]
  assign dot_14_clock = clock; // @[:@18717.4]
  assign dot_14_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19928.4]
  assign dot_14_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19932.4]
  assign dot_14_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19936.4]
  assign dot_14_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19940.4]
  assign dot_14_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19944.4]
  assign dot_14_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19948.4]
  assign dot_14_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19952.4]
  assign dot_14_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19956.4]
  assign dot_14_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19960.4]
  assign dot_14_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19964.4]
  assign dot_14_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19968.4]
  assign dot_14_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19972.4]
  assign dot_14_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19976.4]
  assign dot_14_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19980.4]
  assign dot_14_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19984.4]
  assign dot_14_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19988.4]
  assign dot_14_io_b_0 = $signed(io_wgt_data_bits_14_0); // @[TensorGemm.scala 165:22:@19930.4]
  assign dot_14_io_b_1 = $signed(io_wgt_data_bits_14_1); // @[TensorGemm.scala 165:22:@19934.4]
  assign dot_14_io_b_2 = $signed(io_wgt_data_bits_14_2); // @[TensorGemm.scala 165:22:@19938.4]
  assign dot_14_io_b_3 = $signed(io_wgt_data_bits_14_3); // @[TensorGemm.scala 165:22:@19942.4]
  assign dot_14_io_b_4 = $signed(io_wgt_data_bits_14_4); // @[TensorGemm.scala 165:22:@19946.4]
  assign dot_14_io_b_5 = $signed(io_wgt_data_bits_14_5); // @[TensorGemm.scala 165:22:@19950.4]
  assign dot_14_io_b_6 = $signed(io_wgt_data_bits_14_6); // @[TensorGemm.scala 165:22:@19954.4]
  assign dot_14_io_b_7 = $signed(io_wgt_data_bits_14_7); // @[TensorGemm.scala 165:22:@19958.4]
  assign dot_14_io_b_8 = $signed(io_wgt_data_bits_14_8); // @[TensorGemm.scala 165:22:@19962.4]
  assign dot_14_io_b_9 = $signed(io_wgt_data_bits_14_9); // @[TensorGemm.scala 165:22:@19966.4]
  assign dot_14_io_b_10 = $signed(io_wgt_data_bits_14_10); // @[TensorGemm.scala 165:22:@19970.4]
  assign dot_14_io_b_11 = $signed(io_wgt_data_bits_14_11); // @[TensorGemm.scala 165:22:@19974.4]
  assign dot_14_io_b_12 = $signed(io_wgt_data_bits_14_12); // @[TensorGemm.scala 165:22:@19978.4]
  assign dot_14_io_b_13 = $signed(io_wgt_data_bits_14_13); // @[TensorGemm.scala 165:22:@19982.4]
  assign dot_14_io_b_14 = $signed(io_wgt_data_bits_14_14); // @[TensorGemm.scala 165:22:@19986.4]
  assign dot_14_io_b_15 = $signed(io_wgt_data_bits_14_15); // @[TensorGemm.scala 165:22:@19990.4]
  assign dot_15_clock = clock; // @[:@18720.4]
  assign dot_15_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@20009.4]
  assign dot_15_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@20013.4]
  assign dot_15_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@20017.4]
  assign dot_15_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@20021.4]
  assign dot_15_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@20025.4]
  assign dot_15_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@20029.4]
  assign dot_15_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@20033.4]
  assign dot_15_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@20037.4]
  assign dot_15_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@20041.4]
  assign dot_15_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@20045.4]
  assign dot_15_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@20049.4]
  assign dot_15_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@20053.4]
  assign dot_15_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@20057.4]
  assign dot_15_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@20061.4]
  assign dot_15_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@20065.4]
  assign dot_15_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@20069.4]
  assign dot_15_io_b_0 = $signed(io_wgt_data_bits_15_0); // @[TensorGemm.scala 165:22:@20011.4]
  assign dot_15_io_b_1 = $signed(io_wgt_data_bits_15_1); // @[TensorGemm.scala 165:22:@20015.4]
  assign dot_15_io_b_2 = $signed(io_wgt_data_bits_15_2); // @[TensorGemm.scala 165:22:@20019.4]
  assign dot_15_io_b_3 = $signed(io_wgt_data_bits_15_3); // @[TensorGemm.scala 165:22:@20023.4]
  assign dot_15_io_b_4 = $signed(io_wgt_data_bits_15_4); // @[TensorGemm.scala 165:22:@20027.4]
  assign dot_15_io_b_5 = $signed(io_wgt_data_bits_15_5); // @[TensorGemm.scala 165:22:@20031.4]
  assign dot_15_io_b_6 = $signed(io_wgt_data_bits_15_6); // @[TensorGemm.scala 165:22:@20035.4]
  assign dot_15_io_b_7 = $signed(io_wgt_data_bits_15_7); // @[TensorGemm.scala 165:22:@20039.4]
  assign dot_15_io_b_8 = $signed(io_wgt_data_bits_15_8); // @[TensorGemm.scala 165:22:@20043.4]
  assign dot_15_io_b_9 = $signed(io_wgt_data_bits_15_9); // @[TensorGemm.scala 165:22:@20047.4]
  assign dot_15_io_b_10 = $signed(io_wgt_data_bits_15_10); // @[TensorGemm.scala 165:22:@20051.4]
  assign dot_15_io_b_11 = $signed(io_wgt_data_bits_15_11); // @[TensorGemm.scala 165:22:@20055.4]
  assign dot_15_io_b_12 = $signed(io_wgt_data_bits_15_12); // @[TensorGemm.scala 165:22:@20059.4]
  assign dot_15_io_b_13 = $signed(io_wgt_data_bits_15_13); // @[TensorGemm.scala 165:22:@20063.4]
  assign dot_15_io_b_14 = $signed(io_wgt_data_bits_15_14); // @[TensorGemm.scala 165:22:@20067.4]
  assign dot_15_io_b_15 = $signed(io_wgt_data_bits_15_15); // @[TensorGemm.scala 165:22:@20071.4]
  assign acc_0_clock = clock; // @[:@18723.4]
  assign acc_0_reset = reset; // @[:@18724.4]
  assign acc_0_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@18791.4]
  assign acc_0_io_enq_bits = io_acc_i_data_bits_0_0; // @[TensorGemm.scala 162:24:@18792.4]
  assign acc_1_clock = clock; // @[:@18726.4]
  assign acc_1_reset = reset; // @[:@18727.4]
  assign acc_1_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@18872.4]
  assign acc_1_io_enq_bits = io_acc_i_data_bits_0_1; // @[TensorGemm.scala 162:24:@18873.4]
  assign acc_2_clock = clock; // @[:@18729.4]
  assign acc_2_reset = reset; // @[:@18730.4]
  assign acc_2_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@18953.4]
  assign acc_2_io_enq_bits = io_acc_i_data_bits_0_2; // @[TensorGemm.scala 162:24:@18954.4]
  assign acc_3_clock = clock; // @[:@18732.4]
  assign acc_3_reset = reset; // @[:@18733.4]
  assign acc_3_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19034.4]
  assign acc_3_io_enq_bits = io_acc_i_data_bits_0_3; // @[TensorGemm.scala 162:24:@19035.4]
  assign acc_4_clock = clock; // @[:@18735.4]
  assign acc_4_reset = reset; // @[:@18736.4]
  assign acc_4_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19115.4]
  assign acc_4_io_enq_bits = io_acc_i_data_bits_0_4; // @[TensorGemm.scala 162:24:@19116.4]
  assign acc_5_clock = clock; // @[:@18738.4]
  assign acc_5_reset = reset; // @[:@18739.4]
  assign acc_5_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19196.4]
  assign acc_5_io_enq_bits = io_acc_i_data_bits_0_5; // @[TensorGemm.scala 162:24:@19197.4]
  assign acc_6_clock = clock; // @[:@18741.4]
  assign acc_6_reset = reset; // @[:@18742.4]
  assign acc_6_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19277.4]
  assign acc_6_io_enq_bits = io_acc_i_data_bits_0_6; // @[TensorGemm.scala 162:24:@19278.4]
  assign acc_7_clock = clock; // @[:@18744.4]
  assign acc_7_reset = reset; // @[:@18745.4]
  assign acc_7_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19358.4]
  assign acc_7_io_enq_bits = io_acc_i_data_bits_0_7; // @[TensorGemm.scala 162:24:@19359.4]
  assign acc_8_clock = clock; // @[:@18747.4]
  assign acc_8_reset = reset; // @[:@18748.4]
  assign acc_8_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19439.4]
  assign acc_8_io_enq_bits = io_acc_i_data_bits_0_8; // @[TensorGemm.scala 162:24:@19440.4]
  assign acc_9_clock = clock; // @[:@18750.4]
  assign acc_9_reset = reset; // @[:@18751.4]
  assign acc_9_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19520.4]
  assign acc_9_io_enq_bits = io_acc_i_data_bits_0_9; // @[TensorGemm.scala 162:24:@19521.4]
  assign acc_10_clock = clock; // @[:@18753.4]
  assign acc_10_reset = reset; // @[:@18754.4]
  assign acc_10_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19601.4]
  assign acc_10_io_enq_bits = io_acc_i_data_bits_0_10; // @[TensorGemm.scala 162:24:@19602.4]
  assign acc_11_clock = clock; // @[:@18756.4]
  assign acc_11_reset = reset; // @[:@18757.4]
  assign acc_11_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19682.4]
  assign acc_11_io_enq_bits = io_acc_i_data_bits_0_11; // @[TensorGemm.scala 162:24:@19683.4]
  assign acc_12_clock = clock; // @[:@18759.4]
  assign acc_12_reset = reset; // @[:@18760.4]
  assign acc_12_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19763.4]
  assign acc_12_io_enq_bits = io_acc_i_data_bits_0_12; // @[TensorGemm.scala 162:24:@19764.4]
  assign acc_13_clock = clock; // @[:@18762.4]
  assign acc_13_reset = reset; // @[:@18763.4]
  assign acc_13_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19844.4]
  assign acc_13_io_enq_bits = io_acc_i_data_bits_0_13; // @[TensorGemm.scala 162:24:@19845.4]
  assign acc_14_clock = clock; // @[:@18765.4]
  assign acc_14_reset = reset; // @[:@18766.4]
  assign acc_14_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19925.4]
  assign acc_14_io_enq_bits = io_acc_i_data_bits_0_14; // @[TensorGemm.scala 162:24:@19926.4]
  assign acc_15_clock = clock; // @[:@18768.4]
  assign acc_15_reset = reset; // @[:@18769.4]
  assign acc_15_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@20006.4]
  assign acc_15_io_enq_bits = io_acc_i_data_bits_0_15; // @[TensorGemm.scala 162:24:@20007.4]
endmodule
module Pipe_16( // @[:@20121.2]
  input         clock, // @[:@20122.4]
  input         reset, // @[:@20123.4]
  input         io_enq_valid, // @[:@20124.4]
  input  [13:0] io_enq_bits, // @[:@20124.4]
  output        io_deq_valid, // @[:@20124.4]
  output [13:0] io_deq_bits // @[:@20124.4]
);
  reg  _T_19; // @[Valid.scala 48:22:@20126.4]
  reg [31:0] _RAND_0;
  reg [13:0] _T_21; // @[Reg.scala 11:16:@20128.4]
  reg [31:0] _RAND_1;
  reg  _T_24; // @[Valid.scala 48:22:@20132.4]
  reg [31:0] _RAND_2;
  reg [13:0] _T_26; // @[Reg.scala 11:16:@20134.4]
  reg [31:0] _RAND_3;
  assign io_deq_valid = _T_24; // @[Valid.scala 70:10:@20142.4]
  assign io_deq_bits = _T_26; // @[Valid.scala 70:10:@20141.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_21 = _RAND_1[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_24 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_26 = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      _T_19 <= io_enq_valid;
    end
    if (io_enq_valid) begin
      _T_21 <= io_enq_bits;
    end
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_19;
    end
    if (_T_19) begin
      _T_26 <= _T_21;
    end
  end
endmodule
module TensorGemm( // @[:@20144.2]
  input          clock, // @[:@20145.4]
  input          reset, // @[:@20146.4]
  input          io_start, // @[:@20147.4]
  output         io_done, // @[:@20147.4]
  input  [127:0] io_inst, // @[:@20147.4]
  output         io_uop_idx_valid, // @[:@20147.4]
  output [10:0]  io_uop_idx_bits, // @[:@20147.4]
  input          io_uop_data_valid, // @[:@20147.4]
  input  [9:0]   io_uop_data_bits_u2, // @[:@20147.4]
  input  [10:0]  io_uop_data_bits_u1, // @[:@20147.4]
  input  [10:0]  io_uop_data_bits_u0, // @[:@20147.4]
  output         io_inp_rd_idx_valid, // @[:@20147.4]
  output [10:0]  io_inp_rd_idx_bits, // @[:@20147.4]
  input          io_inp_rd_data_valid, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_0, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_1, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_2, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_3, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_4, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_5, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_6, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_7, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_8, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_9, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_10, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_11, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_12, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_13, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_14, // @[:@20147.4]
  input  [7:0]   io_inp_rd_data_bits_0_15, // @[:@20147.4]
  output         io_wgt_rd_idx_valid, // @[:@20147.4]
  output [9:0]   io_wgt_rd_idx_bits, // @[:@20147.4]
  input          io_wgt_rd_data_valid, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_0_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_1_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_2_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_3_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_4_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_5_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_6_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_7_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_8_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_9_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_10_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_11_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_12_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_13_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_14_15, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_0, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_1, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_2, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_3, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_4, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_5, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_6, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_7, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_8, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_9, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_10, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_11, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_12, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_13, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_14, // @[:@20147.4]
  input  [7:0]   io_wgt_rd_data_bits_15_15, // @[:@20147.4]
  output         io_acc_rd_idx_valid, // @[:@20147.4]
  output [10:0]  io_acc_rd_idx_bits, // @[:@20147.4]
  input          io_acc_rd_data_valid, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_0, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_1, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_2, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_3, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_4, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_5, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_6, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_7, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_8, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_9, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_10, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_11, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_12, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_13, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_14, // @[:@20147.4]
  input  [31:0]  io_acc_rd_data_bits_0_15, // @[:@20147.4]
  output         io_acc_wr_valid, // @[:@20147.4]
  output [10:0]  io_acc_wr_bits_idx, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_0, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_1, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_2, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_3, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_4, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_5, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_6, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_7, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_8, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_9, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_10, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_11, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_12, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_13, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_14, // @[:@20147.4]
  output [31:0]  io_acc_wr_bits_data_0_15, // @[:@20147.4]
  output         io_out_wr_valid, // @[:@20147.4]
  output [10:0]  io_out_wr_bits_idx, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_0, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_1, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_2, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_3, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_4, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_5, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_6, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_7, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_8, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_9, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_10, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_11, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_12, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_13, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_14, // @[:@20147.4]
  output [7:0]   io_out_wr_bits_data_0_15 // @[:@20147.4]
);
  wire  mvc_clock; // @[TensorGemm.scala 199:19:@20150.4]
  wire  mvc_reset; // @[TensorGemm.scala 199:19:@20150.4]
  wire  mvc_io_reset; // @[TensorGemm.scala 199:19:@20150.4]
  wire  mvc_io_inp_data_valid; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_inp_data_bits_0_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire  mvc_io_wgt_data_valid; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_0_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_1_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_2_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_3_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_4_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_5_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_6_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_7_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_8_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_9_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_10_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_11_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_12_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_13_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_14_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_wgt_data_bits_15_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire  mvc_io_acc_i_data_valid; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire  mvc_io_acc_o_data_valid; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire  mvc_io_out_data_valid; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_0; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_1; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_2; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_3; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_4; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_5; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_6; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_7; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_8; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_9; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_10; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_11; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_12; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_13; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_14; // @[TensorGemm.scala 199:19:@20150.4]
  wire [7:0] mvc_io_out_data_bits_0_15; // @[TensorGemm.scala 199:19:@20150.4]
  wire  wrpipe_clock; // @[TensorGemm.scala 218:22:@20203.4]
  wire  wrpipe_reset; // @[TensorGemm.scala 218:22:@20203.4]
  wire  wrpipe_io_enq_valid; // @[TensorGemm.scala 218:22:@20203.4]
  wire [13:0] wrpipe_io_enq_bits; // @[TensorGemm.scala 218:22:@20203.4]
  wire  wrpipe_io_deq_valid; // @[TensorGemm.scala 218:22:@20203.4]
  wire [13:0] wrpipe_io_deq_bits; // @[TensorGemm.scala 218:22:@20203.4]
  reg [2:0] state; // @[TensorGemm.scala 198:22:@20149.4]
  reg [31:0] _RAND_0;
  wire  dec_reset; // @[TensorGemm.scala 200:29:@20166.4]
  wire [12:0] dec_uop_begin; // @[TensorGemm.scala 200:29:@20168.4]
  wire [13:0] dec_uop_end; // @[TensorGemm.scala 200:29:@20170.4]
  wire [13:0] dec_lp_0; // @[TensorGemm.scala 200:29:@20172.4]
  wire [13:0] dec_lp_1; // @[TensorGemm.scala 200:29:@20174.4]
  wire [10:0] dec_acc_0; // @[TensorGemm.scala 200:29:@20178.4]
  wire [10:0] dec_acc_1; // @[TensorGemm.scala 200:29:@20180.4]
  wire [10:0] dec_inp_0; // @[TensorGemm.scala 200:29:@20182.4]
  wire [10:0] dec_inp_1; // @[TensorGemm.scala 200:29:@20184.4]
  wire [9:0] dec_wgt_0; // @[TensorGemm.scala 200:29:@20186.4]
  wire [9:0] dec_wgt_1; // @[TensorGemm.scala 200:29:@20188.4]
  reg [13:0] uop_idx; // @[TensorGemm.scala 201:20:@20190.4]
  reg [31:0] _RAND_1;
  reg [13:0] uop_acc; // @[TensorGemm.scala 203:20:@20191.4]
  reg [31:0] _RAND_2;
  reg [13:0] uop_inp; // @[TensorGemm.scala 204:20:@20192.4]
  reg [31:0] _RAND_3;
  reg [13:0] uop_wgt; // @[TensorGemm.scala 205:20:@20193.4]
  reg [31:0] _RAND_4;
  reg [13:0] cnt_o; // @[TensorGemm.scala 206:18:@20194.4]
  reg [31:0] _RAND_5;
  reg [13:0] acc_o; // @[TensorGemm.scala 207:18:@20195.4]
  reg [31:0] _RAND_6;
  reg [13:0] inp_o; // @[TensorGemm.scala 208:18:@20196.4]
  reg [31:0] _RAND_7;
  reg [13:0] wgt_o; // @[TensorGemm.scala 209:18:@20197.4]
  reg [31:0] _RAND_8;
  reg [13:0] cnt_i; // @[TensorGemm.scala 210:18:@20198.4]
  reg [31:0] _RAND_9;
  reg [13:0] acc_i; // @[TensorGemm.scala 211:18:@20199.4]
  reg [31:0] _RAND_10;
  reg [13:0] inp_i; // @[TensorGemm.scala 212:18:@20200.4]
  reg [31:0] _RAND_11;
  reg [13:0] wgt_i; // @[TensorGemm.scala 213:18:@20201.4]
  reg [31:0] _RAND_12;
  reg [4:0] inflight; // @[TensorGemm.scala 215:21:@20202.4]
  reg [31:0] _RAND_13;
  wire  _T_7688; // @[TensorGemm.scala 219:23:@20206.4]
  wire  _T_7689; // @[TensorGemm.scala 220:13:@20207.4]
  wire [14:0] _T_7691; // @[TensorGemm.scala 221:26:@20208.4]
  wire [14:0] _T_7692; // @[TensorGemm.scala 221:26:@20209.4]
  wire [13:0] _T_7693; // @[TensorGemm.scala 221:26:@20210.4]
  wire  _T_7694; // @[TensorGemm.scala 221:13:@20211.4]
  wire  _T_7695; // @[TensorGemm.scala 220:22:@20212.4]
  wire [14:0] _T_7697; // @[TensorGemm.scala 222:26:@20213.4]
  wire [14:0] _T_7698; // @[TensorGemm.scala 222:26:@20214.4]
  wire [13:0] _T_7699; // @[TensorGemm.scala 222:26:@20215.4]
  wire  _T_7700; // @[TensorGemm.scala 222:13:@20216.4]
  wire  _T_7701; // @[TensorGemm.scala 221:32:@20217.4]
  wire [14:0] _T_7703; // @[TensorGemm.scala 223:27:@20218.4]
  wire [14:0] _T_7704; // @[TensorGemm.scala 223:27:@20219.4]
  wire [13:0] _T_7705; // @[TensorGemm.scala 223:27:@20220.4]
  wire  _T_7706; // @[TensorGemm.scala 223:15:@20221.4]
  wire  _T_7707; // @[TensorGemm.scala 222:32:@20222.4]
  wire  _T_7710; // @[TensorGemm.scala 223:33:@20224.4]
  wire  _T_7711; // @[TensorGemm.scala 225:13:@20225.4]
  wire  _T_7712; // @[TensorGemm.scala 224:25:@20226.4]
  wire  _T_7713; // @[Conditional.scala 37:30:@20228.4]
  wire [2:0] _GEN_0; // @[TensorGemm.scala 229:22:@20230.6]
  wire  _T_7714; // @[Conditional.scala 37:30:@20235.6]
  wire  _T_7715; // @[Conditional.scala 37:30:@20240.8]
  wire  _T_7716; // @[Conditional.scala 37:30:@20245.10]
  wire  _T_7717; // @[Conditional.scala 37:30:@20250.12]
  wire  _T_7728; // @[TensorGemm.scala 244:36:@20260.14]
  wire  _T_7734; // @[TensorGemm.scala 245:38:@20265.14]
  wire  _T_7736; // @[TensorGemm.scala 247:23:@20267.16]
  wire [2:0] _GEN_1; // @[TensorGemm.scala 247:32:@20268.16]
  wire [2:0] _GEN_2; // @[TensorGemm.scala 246:40:@20266.14]
  wire  _T_7737; // @[Conditional.scala 37:30:@20280.14]
  wire [2:0] _GEN_3; // @[TensorGemm.scala 257:30:@20283.16]
  wire [2:0] _GEN_4; // @[Conditional.scala 39:67:@20281.14]
  wire [2:0] _GEN_5; // @[Conditional.scala 39:67:@20251.12]
  wire [2:0] _GEN_6; // @[Conditional.scala 39:67:@20246.10]
  wire [2:0] _GEN_7; // @[Conditional.scala 39:67:@20241.8]
  wire [2:0] _GEN_8; // @[Conditional.scala 39:67:@20236.6]
  wire [2:0] _GEN_9; // @[Conditional.scala 40:58:@20229.4]
  wire  _T_7740; // @[TensorGemm.scala 263:14:@20287.4]
  wire  _T_7743; // @[TensorGemm.scala 265:14:@20292.6]
  wire  _T_7744; // @[TensorGemm.scala 266:17:@20294.8]
  wire  _T_7745; // @[TensorGemm.scala 266:34:@20295.8]
  wire [5:0] _T_7748; // @[TensorGemm.scala 269:28:@20302.12]
  wire [4:0] _T_7749; // @[TensorGemm.scala 269:28:@20303.12]
  wire [5:0] _T_7751; // @[TensorGemm.scala 271:28:@20308.14]
  wire [5:0] _T_7752; // @[TensorGemm.scala 271:28:@20309.14]
  wire [4:0] _T_7753; // @[TensorGemm.scala 271:28:@20310.14]
  wire [4:0] _GEN_10; // @[TensorGemm.scala 270:41:@20307.12]
  wire [4:0] _GEN_11; // @[TensorGemm.scala 268:39:@20301.10]
  wire [4:0] _GEN_12; // @[TensorGemm.scala 266:62:@20296.8]
  wire [4:0] _GEN_13; // @[TensorGemm.scala 265:26:@20293.6]
  wire  _T_7761; // @[TensorGemm.scala 277:23:@20320.4]
  wire  _T_7762; // @[TensorGemm.scala 276:21:@20321.4]
  wire [13:0] _GEN_40; // @[TensorGemm.scala 280:46:@20327.6]
  wire  _T_7764; // @[TensorGemm.scala 280:46:@20327.6]
  wire  _T_7765; // @[TensorGemm.scala 280:29:@20328.6]
  wire [14:0] _T_7767; // @[TensorGemm.scala 281:24:@20330.8]
  wire [13:0] _T_7768; // @[TensorGemm.scala 281:24:@20331.8]
  wire [13:0] _GEN_15; // @[TensorGemm.scala 280:59:@20329.6]
  wire  _T_7786; // @[TensorGemm.scala 291:33:@20352.6]
  wire [14:0] _T_7788; // @[TensorGemm.scala 293:20:@20354.8]
  wire [13:0] _T_7789; // @[TensorGemm.scala 293:20:@20355.8]
  wire [13:0] _GEN_41; // @[TensorGemm.scala 294:20:@20357.8]
  wire [14:0] _T_7790; // @[TensorGemm.scala 294:20:@20357.8]
  wire [13:0] _T_7791; // @[TensorGemm.scala 294:20:@20358.8]
  wire [13:0] _GEN_42; // @[TensorGemm.scala 295:20:@20360.8]
  wire [14:0] _T_7792; // @[TensorGemm.scala 295:20:@20360.8]
  wire [13:0] _T_7793; // @[TensorGemm.scala 295:20:@20361.8]
  wire [13:0] _GEN_43; // @[TensorGemm.scala 296:20:@20363.8]
  wire [14:0] _T_7794; // @[TensorGemm.scala 296:20:@20363.8]
  wire [13:0] _T_7795; // @[TensorGemm.scala 296:20:@20364.8]
  wire [13:0] _GEN_17; // @[TensorGemm.scala 292:33:@20353.6]
  wire [13:0] _GEN_18; // @[TensorGemm.scala 292:33:@20353.6]
  wire [13:0] _GEN_19; // @[TensorGemm.scala 292:33:@20353.6]
  wire [13:0] _GEN_20; // @[TensorGemm.scala 292:33:@20353.6]
  wire  _T_7801; // @[TensorGemm.scala 304:20:@20375.6]
  wire  _T_7802; // @[TensorGemm.scala 304:42:@20376.6]
  wire  _T_7803; // @[TensorGemm.scala 304:33:@20377.6]
  wire [14:0] _T_7813; // @[TensorGemm.scala 310:20:@20392.10]
  wire [13:0] _T_7814; // @[TensorGemm.scala 310:20:@20393.10]
  wire [13:0] _GEN_44; // @[TensorGemm.scala 311:20:@20395.10]
  wire [14:0] _T_7815; // @[TensorGemm.scala 311:20:@20395.10]
  wire [13:0] _T_7816; // @[TensorGemm.scala 311:20:@20396.10]
  wire [13:0] _GEN_45; // @[TensorGemm.scala 312:20:@20398.10]
  wire [14:0] _T_7817; // @[TensorGemm.scala 312:20:@20398.10]
  wire [13:0] _T_7818; // @[TensorGemm.scala 312:20:@20399.10]
  wire [13:0] _GEN_46; // @[TensorGemm.scala 313:20:@20401.10]
  wire [14:0] _T_7819; // @[TensorGemm.scala 313:20:@20401.10]
  wire [13:0] _T_7820; // @[TensorGemm.scala 313:20:@20402.10]
  wire [13:0] _GEN_25; // @[TensorGemm.scala 309:59:@20391.8]
  wire [13:0] _GEN_26; // @[TensorGemm.scala 309:59:@20391.8]
  wire [13:0] _GEN_27; // @[TensorGemm.scala 309:59:@20391.8]
  wire [13:0] _GEN_28; // @[TensorGemm.scala 309:59:@20391.8]
  wire [13:0] _GEN_29; // @[TensorGemm.scala 304:56:@20378.6]
  wire [13:0] _GEN_30; // @[TensorGemm.scala 304:56:@20378.6]
  wire [13:0] _GEN_31; // @[TensorGemm.scala 304:56:@20378.6]
  wire [13:0] _GEN_32; // @[TensorGemm.scala 304:56:@20378.6]
  wire  _T_7821; // @[TensorGemm.scala 316:14:@20405.4]
  wire  _T_7822; // @[TensorGemm.scala 316:30:@20406.4]
  wire [13:0] _GEN_47; // @[TensorGemm.scala 317:36:@20408.6]
  wire [14:0] _T_7823; // @[TensorGemm.scala 317:36:@20408.6]
  wire [13:0] _T_7824; // @[TensorGemm.scala 317:36:@20409.6]
  wire [13:0] _GEN_48; // @[TensorGemm.scala 318:36:@20411.6]
  wire [14:0] _T_7825; // @[TensorGemm.scala 318:36:@20411.6]
  wire [13:0] _T_7826; // @[TensorGemm.scala 318:36:@20412.6]
  wire [13:0] _GEN_49; // @[TensorGemm.scala 319:36:@20414.6]
  wire [14:0] _T_7827; // @[TensorGemm.scala 319:36:@20414.6]
  wire [13:0] _T_7828; // @[TensorGemm.scala 319:36:@20415.6]
  wire  _T_7830; // @[TensorGemm.scala 322:43:@20419.4]
  wire  _T_8115; // @[TensorGemm.scala 351:8:@21005.4]
  wire [13:0] _T_8117; // @[TensorGemm.scala 352:28:@21008.4]
  MatrixVectorMultiplication mvc ( // @[TensorGemm.scala 199:19:@20150.4]
    .clock(mvc_clock),
    .reset(mvc_reset),
    .io_reset(mvc_io_reset),
    .io_inp_data_valid(mvc_io_inp_data_valid),
    .io_inp_data_bits_0_0(mvc_io_inp_data_bits_0_0),
    .io_inp_data_bits_0_1(mvc_io_inp_data_bits_0_1),
    .io_inp_data_bits_0_2(mvc_io_inp_data_bits_0_2),
    .io_inp_data_bits_0_3(mvc_io_inp_data_bits_0_3),
    .io_inp_data_bits_0_4(mvc_io_inp_data_bits_0_4),
    .io_inp_data_bits_0_5(mvc_io_inp_data_bits_0_5),
    .io_inp_data_bits_0_6(mvc_io_inp_data_bits_0_6),
    .io_inp_data_bits_0_7(mvc_io_inp_data_bits_0_7),
    .io_inp_data_bits_0_8(mvc_io_inp_data_bits_0_8),
    .io_inp_data_bits_0_9(mvc_io_inp_data_bits_0_9),
    .io_inp_data_bits_0_10(mvc_io_inp_data_bits_0_10),
    .io_inp_data_bits_0_11(mvc_io_inp_data_bits_0_11),
    .io_inp_data_bits_0_12(mvc_io_inp_data_bits_0_12),
    .io_inp_data_bits_0_13(mvc_io_inp_data_bits_0_13),
    .io_inp_data_bits_0_14(mvc_io_inp_data_bits_0_14),
    .io_inp_data_bits_0_15(mvc_io_inp_data_bits_0_15),
    .io_wgt_data_valid(mvc_io_wgt_data_valid),
    .io_wgt_data_bits_0_0(mvc_io_wgt_data_bits_0_0),
    .io_wgt_data_bits_0_1(mvc_io_wgt_data_bits_0_1),
    .io_wgt_data_bits_0_2(mvc_io_wgt_data_bits_0_2),
    .io_wgt_data_bits_0_3(mvc_io_wgt_data_bits_0_3),
    .io_wgt_data_bits_0_4(mvc_io_wgt_data_bits_0_4),
    .io_wgt_data_bits_0_5(mvc_io_wgt_data_bits_0_5),
    .io_wgt_data_bits_0_6(mvc_io_wgt_data_bits_0_6),
    .io_wgt_data_bits_0_7(mvc_io_wgt_data_bits_0_7),
    .io_wgt_data_bits_0_8(mvc_io_wgt_data_bits_0_8),
    .io_wgt_data_bits_0_9(mvc_io_wgt_data_bits_0_9),
    .io_wgt_data_bits_0_10(mvc_io_wgt_data_bits_0_10),
    .io_wgt_data_bits_0_11(mvc_io_wgt_data_bits_0_11),
    .io_wgt_data_bits_0_12(mvc_io_wgt_data_bits_0_12),
    .io_wgt_data_bits_0_13(mvc_io_wgt_data_bits_0_13),
    .io_wgt_data_bits_0_14(mvc_io_wgt_data_bits_0_14),
    .io_wgt_data_bits_0_15(mvc_io_wgt_data_bits_0_15),
    .io_wgt_data_bits_1_0(mvc_io_wgt_data_bits_1_0),
    .io_wgt_data_bits_1_1(mvc_io_wgt_data_bits_1_1),
    .io_wgt_data_bits_1_2(mvc_io_wgt_data_bits_1_2),
    .io_wgt_data_bits_1_3(mvc_io_wgt_data_bits_1_3),
    .io_wgt_data_bits_1_4(mvc_io_wgt_data_bits_1_4),
    .io_wgt_data_bits_1_5(mvc_io_wgt_data_bits_1_5),
    .io_wgt_data_bits_1_6(mvc_io_wgt_data_bits_1_6),
    .io_wgt_data_bits_1_7(mvc_io_wgt_data_bits_1_7),
    .io_wgt_data_bits_1_8(mvc_io_wgt_data_bits_1_8),
    .io_wgt_data_bits_1_9(mvc_io_wgt_data_bits_1_9),
    .io_wgt_data_bits_1_10(mvc_io_wgt_data_bits_1_10),
    .io_wgt_data_bits_1_11(mvc_io_wgt_data_bits_1_11),
    .io_wgt_data_bits_1_12(mvc_io_wgt_data_bits_1_12),
    .io_wgt_data_bits_1_13(mvc_io_wgt_data_bits_1_13),
    .io_wgt_data_bits_1_14(mvc_io_wgt_data_bits_1_14),
    .io_wgt_data_bits_1_15(mvc_io_wgt_data_bits_1_15),
    .io_wgt_data_bits_2_0(mvc_io_wgt_data_bits_2_0),
    .io_wgt_data_bits_2_1(mvc_io_wgt_data_bits_2_1),
    .io_wgt_data_bits_2_2(mvc_io_wgt_data_bits_2_2),
    .io_wgt_data_bits_2_3(mvc_io_wgt_data_bits_2_3),
    .io_wgt_data_bits_2_4(mvc_io_wgt_data_bits_2_4),
    .io_wgt_data_bits_2_5(mvc_io_wgt_data_bits_2_5),
    .io_wgt_data_bits_2_6(mvc_io_wgt_data_bits_2_6),
    .io_wgt_data_bits_2_7(mvc_io_wgt_data_bits_2_7),
    .io_wgt_data_bits_2_8(mvc_io_wgt_data_bits_2_8),
    .io_wgt_data_bits_2_9(mvc_io_wgt_data_bits_2_9),
    .io_wgt_data_bits_2_10(mvc_io_wgt_data_bits_2_10),
    .io_wgt_data_bits_2_11(mvc_io_wgt_data_bits_2_11),
    .io_wgt_data_bits_2_12(mvc_io_wgt_data_bits_2_12),
    .io_wgt_data_bits_2_13(mvc_io_wgt_data_bits_2_13),
    .io_wgt_data_bits_2_14(mvc_io_wgt_data_bits_2_14),
    .io_wgt_data_bits_2_15(mvc_io_wgt_data_bits_2_15),
    .io_wgt_data_bits_3_0(mvc_io_wgt_data_bits_3_0),
    .io_wgt_data_bits_3_1(mvc_io_wgt_data_bits_3_1),
    .io_wgt_data_bits_3_2(mvc_io_wgt_data_bits_3_2),
    .io_wgt_data_bits_3_3(mvc_io_wgt_data_bits_3_3),
    .io_wgt_data_bits_3_4(mvc_io_wgt_data_bits_3_4),
    .io_wgt_data_bits_3_5(mvc_io_wgt_data_bits_3_5),
    .io_wgt_data_bits_3_6(mvc_io_wgt_data_bits_3_6),
    .io_wgt_data_bits_3_7(mvc_io_wgt_data_bits_3_7),
    .io_wgt_data_bits_3_8(mvc_io_wgt_data_bits_3_8),
    .io_wgt_data_bits_3_9(mvc_io_wgt_data_bits_3_9),
    .io_wgt_data_bits_3_10(mvc_io_wgt_data_bits_3_10),
    .io_wgt_data_bits_3_11(mvc_io_wgt_data_bits_3_11),
    .io_wgt_data_bits_3_12(mvc_io_wgt_data_bits_3_12),
    .io_wgt_data_bits_3_13(mvc_io_wgt_data_bits_3_13),
    .io_wgt_data_bits_3_14(mvc_io_wgt_data_bits_3_14),
    .io_wgt_data_bits_3_15(mvc_io_wgt_data_bits_3_15),
    .io_wgt_data_bits_4_0(mvc_io_wgt_data_bits_4_0),
    .io_wgt_data_bits_4_1(mvc_io_wgt_data_bits_4_1),
    .io_wgt_data_bits_4_2(mvc_io_wgt_data_bits_4_2),
    .io_wgt_data_bits_4_3(mvc_io_wgt_data_bits_4_3),
    .io_wgt_data_bits_4_4(mvc_io_wgt_data_bits_4_4),
    .io_wgt_data_bits_4_5(mvc_io_wgt_data_bits_4_5),
    .io_wgt_data_bits_4_6(mvc_io_wgt_data_bits_4_6),
    .io_wgt_data_bits_4_7(mvc_io_wgt_data_bits_4_7),
    .io_wgt_data_bits_4_8(mvc_io_wgt_data_bits_4_8),
    .io_wgt_data_bits_4_9(mvc_io_wgt_data_bits_4_9),
    .io_wgt_data_bits_4_10(mvc_io_wgt_data_bits_4_10),
    .io_wgt_data_bits_4_11(mvc_io_wgt_data_bits_4_11),
    .io_wgt_data_bits_4_12(mvc_io_wgt_data_bits_4_12),
    .io_wgt_data_bits_4_13(mvc_io_wgt_data_bits_4_13),
    .io_wgt_data_bits_4_14(mvc_io_wgt_data_bits_4_14),
    .io_wgt_data_bits_4_15(mvc_io_wgt_data_bits_4_15),
    .io_wgt_data_bits_5_0(mvc_io_wgt_data_bits_5_0),
    .io_wgt_data_bits_5_1(mvc_io_wgt_data_bits_5_1),
    .io_wgt_data_bits_5_2(mvc_io_wgt_data_bits_5_2),
    .io_wgt_data_bits_5_3(mvc_io_wgt_data_bits_5_3),
    .io_wgt_data_bits_5_4(mvc_io_wgt_data_bits_5_4),
    .io_wgt_data_bits_5_5(mvc_io_wgt_data_bits_5_5),
    .io_wgt_data_bits_5_6(mvc_io_wgt_data_bits_5_6),
    .io_wgt_data_bits_5_7(mvc_io_wgt_data_bits_5_7),
    .io_wgt_data_bits_5_8(mvc_io_wgt_data_bits_5_8),
    .io_wgt_data_bits_5_9(mvc_io_wgt_data_bits_5_9),
    .io_wgt_data_bits_5_10(mvc_io_wgt_data_bits_5_10),
    .io_wgt_data_bits_5_11(mvc_io_wgt_data_bits_5_11),
    .io_wgt_data_bits_5_12(mvc_io_wgt_data_bits_5_12),
    .io_wgt_data_bits_5_13(mvc_io_wgt_data_bits_5_13),
    .io_wgt_data_bits_5_14(mvc_io_wgt_data_bits_5_14),
    .io_wgt_data_bits_5_15(mvc_io_wgt_data_bits_5_15),
    .io_wgt_data_bits_6_0(mvc_io_wgt_data_bits_6_0),
    .io_wgt_data_bits_6_1(mvc_io_wgt_data_bits_6_1),
    .io_wgt_data_bits_6_2(mvc_io_wgt_data_bits_6_2),
    .io_wgt_data_bits_6_3(mvc_io_wgt_data_bits_6_3),
    .io_wgt_data_bits_6_4(mvc_io_wgt_data_bits_6_4),
    .io_wgt_data_bits_6_5(mvc_io_wgt_data_bits_6_5),
    .io_wgt_data_bits_6_6(mvc_io_wgt_data_bits_6_6),
    .io_wgt_data_bits_6_7(mvc_io_wgt_data_bits_6_7),
    .io_wgt_data_bits_6_8(mvc_io_wgt_data_bits_6_8),
    .io_wgt_data_bits_6_9(mvc_io_wgt_data_bits_6_9),
    .io_wgt_data_bits_6_10(mvc_io_wgt_data_bits_6_10),
    .io_wgt_data_bits_6_11(mvc_io_wgt_data_bits_6_11),
    .io_wgt_data_bits_6_12(mvc_io_wgt_data_bits_6_12),
    .io_wgt_data_bits_6_13(mvc_io_wgt_data_bits_6_13),
    .io_wgt_data_bits_6_14(mvc_io_wgt_data_bits_6_14),
    .io_wgt_data_bits_6_15(mvc_io_wgt_data_bits_6_15),
    .io_wgt_data_bits_7_0(mvc_io_wgt_data_bits_7_0),
    .io_wgt_data_bits_7_1(mvc_io_wgt_data_bits_7_1),
    .io_wgt_data_bits_7_2(mvc_io_wgt_data_bits_7_2),
    .io_wgt_data_bits_7_3(mvc_io_wgt_data_bits_7_3),
    .io_wgt_data_bits_7_4(mvc_io_wgt_data_bits_7_4),
    .io_wgt_data_bits_7_5(mvc_io_wgt_data_bits_7_5),
    .io_wgt_data_bits_7_6(mvc_io_wgt_data_bits_7_6),
    .io_wgt_data_bits_7_7(mvc_io_wgt_data_bits_7_7),
    .io_wgt_data_bits_7_8(mvc_io_wgt_data_bits_7_8),
    .io_wgt_data_bits_7_9(mvc_io_wgt_data_bits_7_9),
    .io_wgt_data_bits_7_10(mvc_io_wgt_data_bits_7_10),
    .io_wgt_data_bits_7_11(mvc_io_wgt_data_bits_7_11),
    .io_wgt_data_bits_7_12(mvc_io_wgt_data_bits_7_12),
    .io_wgt_data_bits_7_13(mvc_io_wgt_data_bits_7_13),
    .io_wgt_data_bits_7_14(mvc_io_wgt_data_bits_7_14),
    .io_wgt_data_bits_7_15(mvc_io_wgt_data_bits_7_15),
    .io_wgt_data_bits_8_0(mvc_io_wgt_data_bits_8_0),
    .io_wgt_data_bits_8_1(mvc_io_wgt_data_bits_8_1),
    .io_wgt_data_bits_8_2(mvc_io_wgt_data_bits_8_2),
    .io_wgt_data_bits_8_3(mvc_io_wgt_data_bits_8_3),
    .io_wgt_data_bits_8_4(mvc_io_wgt_data_bits_8_4),
    .io_wgt_data_bits_8_5(mvc_io_wgt_data_bits_8_5),
    .io_wgt_data_bits_8_6(mvc_io_wgt_data_bits_8_6),
    .io_wgt_data_bits_8_7(mvc_io_wgt_data_bits_8_7),
    .io_wgt_data_bits_8_8(mvc_io_wgt_data_bits_8_8),
    .io_wgt_data_bits_8_9(mvc_io_wgt_data_bits_8_9),
    .io_wgt_data_bits_8_10(mvc_io_wgt_data_bits_8_10),
    .io_wgt_data_bits_8_11(mvc_io_wgt_data_bits_8_11),
    .io_wgt_data_bits_8_12(mvc_io_wgt_data_bits_8_12),
    .io_wgt_data_bits_8_13(mvc_io_wgt_data_bits_8_13),
    .io_wgt_data_bits_8_14(mvc_io_wgt_data_bits_8_14),
    .io_wgt_data_bits_8_15(mvc_io_wgt_data_bits_8_15),
    .io_wgt_data_bits_9_0(mvc_io_wgt_data_bits_9_0),
    .io_wgt_data_bits_9_1(mvc_io_wgt_data_bits_9_1),
    .io_wgt_data_bits_9_2(mvc_io_wgt_data_bits_9_2),
    .io_wgt_data_bits_9_3(mvc_io_wgt_data_bits_9_3),
    .io_wgt_data_bits_9_4(mvc_io_wgt_data_bits_9_4),
    .io_wgt_data_bits_9_5(mvc_io_wgt_data_bits_9_5),
    .io_wgt_data_bits_9_6(mvc_io_wgt_data_bits_9_6),
    .io_wgt_data_bits_9_7(mvc_io_wgt_data_bits_9_7),
    .io_wgt_data_bits_9_8(mvc_io_wgt_data_bits_9_8),
    .io_wgt_data_bits_9_9(mvc_io_wgt_data_bits_9_9),
    .io_wgt_data_bits_9_10(mvc_io_wgt_data_bits_9_10),
    .io_wgt_data_bits_9_11(mvc_io_wgt_data_bits_9_11),
    .io_wgt_data_bits_9_12(mvc_io_wgt_data_bits_9_12),
    .io_wgt_data_bits_9_13(mvc_io_wgt_data_bits_9_13),
    .io_wgt_data_bits_9_14(mvc_io_wgt_data_bits_9_14),
    .io_wgt_data_bits_9_15(mvc_io_wgt_data_bits_9_15),
    .io_wgt_data_bits_10_0(mvc_io_wgt_data_bits_10_0),
    .io_wgt_data_bits_10_1(mvc_io_wgt_data_bits_10_1),
    .io_wgt_data_bits_10_2(mvc_io_wgt_data_bits_10_2),
    .io_wgt_data_bits_10_3(mvc_io_wgt_data_bits_10_3),
    .io_wgt_data_bits_10_4(mvc_io_wgt_data_bits_10_4),
    .io_wgt_data_bits_10_5(mvc_io_wgt_data_bits_10_5),
    .io_wgt_data_bits_10_6(mvc_io_wgt_data_bits_10_6),
    .io_wgt_data_bits_10_7(mvc_io_wgt_data_bits_10_7),
    .io_wgt_data_bits_10_8(mvc_io_wgt_data_bits_10_8),
    .io_wgt_data_bits_10_9(mvc_io_wgt_data_bits_10_9),
    .io_wgt_data_bits_10_10(mvc_io_wgt_data_bits_10_10),
    .io_wgt_data_bits_10_11(mvc_io_wgt_data_bits_10_11),
    .io_wgt_data_bits_10_12(mvc_io_wgt_data_bits_10_12),
    .io_wgt_data_bits_10_13(mvc_io_wgt_data_bits_10_13),
    .io_wgt_data_bits_10_14(mvc_io_wgt_data_bits_10_14),
    .io_wgt_data_bits_10_15(mvc_io_wgt_data_bits_10_15),
    .io_wgt_data_bits_11_0(mvc_io_wgt_data_bits_11_0),
    .io_wgt_data_bits_11_1(mvc_io_wgt_data_bits_11_1),
    .io_wgt_data_bits_11_2(mvc_io_wgt_data_bits_11_2),
    .io_wgt_data_bits_11_3(mvc_io_wgt_data_bits_11_3),
    .io_wgt_data_bits_11_4(mvc_io_wgt_data_bits_11_4),
    .io_wgt_data_bits_11_5(mvc_io_wgt_data_bits_11_5),
    .io_wgt_data_bits_11_6(mvc_io_wgt_data_bits_11_6),
    .io_wgt_data_bits_11_7(mvc_io_wgt_data_bits_11_7),
    .io_wgt_data_bits_11_8(mvc_io_wgt_data_bits_11_8),
    .io_wgt_data_bits_11_9(mvc_io_wgt_data_bits_11_9),
    .io_wgt_data_bits_11_10(mvc_io_wgt_data_bits_11_10),
    .io_wgt_data_bits_11_11(mvc_io_wgt_data_bits_11_11),
    .io_wgt_data_bits_11_12(mvc_io_wgt_data_bits_11_12),
    .io_wgt_data_bits_11_13(mvc_io_wgt_data_bits_11_13),
    .io_wgt_data_bits_11_14(mvc_io_wgt_data_bits_11_14),
    .io_wgt_data_bits_11_15(mvc_io_wgt_data_bits_11_15),
    .io_wgt_data_bits_12_0(mvc_io_wgt_data_bits_12_0),
    .io_wgt_data_bits_12_1(mvc_io_wgt_data_bits_12_1),
    .io_wgt_data_bits_12_2(mvc_io_wgt_data_bits_12_2),
    .io_wgt_data_bits_12_3(mvc_io_wgt_data_bits_12_3),
    .io_wgt_data_bits_12_4(mvc_io_wgt_data_bits_12_4),
    .io_wgt_data_bits_12_5(mvc_io_wgt_data_bits_12_5),
    .io_wgt_data_bits_12_6(mvc_io_wgt_data_bits_12_6),
    .io_wgt_data_bits_12_7(mvc_io_wgt_data_bits_12_7),
    .io_wgt_data_bits_12_8(mvc_io_wgt_data_bits_12_8),
    .io_wgt_data_bits_12_9(mvc_io_wgt_data_bits_12_9),
    .io_wgt_data_bits_12_10(mvc_io_wgt_data_bits_12_10),
    .io_wgt_data_bits_12_11(mvc_io_wgt_data_bits_12_11),
    .io_wgt_data_bits_12_12(mvc_io_wgt_data_bits_12_12),
    .io_wgt_data_bits_12_13(mvc_io_wgt_data_bits_12_13),
    .io_wgt_data_bits_12_14(mvc_io_wgt_data_bits_12_14),
    .io_wgt_data_bits_12_15(mvc_io_wgt_data_bits_12_15),
    .io_wgt_data_bits_13_0(mvc_io_wgt_data_bits_13_0),
    .io_wgt_data_bits_13_1(mvc_io_wgt_data_bits_13_1),
    .io_wgt_data_bits_13_2(mvc_io_wgt_data_bits_13_2),
    .io_wgt_data_bits_13_3(mvc_io_wgt_data_bits_13_3),
    .io_wgt_data_bits_13_4(mvc_io_wgt_data_bits_13_4),
    .io_wgt_data_bits_13_5(mvc_io_wgt_data_bits_13_5),
    .io_wgt_data_bits_13_6(mvc_io_wgt_data_bits_13_6),
    .io_wgt_data_bits_13_7(mvc_io_wgt_data_bits_13_7),
    .io_wgt_data_bits_13_8(mvc_io_wgt_data_bits_13_8),
    .io_wgt_data_bits_13_9(mvc_io_wgt_data_bits_13_9),
    .io_wgt_data_bits_13_10(mvc_io_wgt_data_bits_13_10),
    .io_wgt_data_bits_13_11(mvc_io_wgt_data_bits_13_11),
    .io_wgt_data_bits_13_12(mvc_io_wgt_data_bits_13_12),
    .io_wgt_data_bits_13_13(mvc_io_wgt_data_bits_13_13),
    .io_wgt_data_bits_13_14(mvc_io_wgt_data_bits_13_14),
    .io_wgt_data_bits_13_15(mvc_io_wgt_data_bits_13_15),
    .io_wgt_data_bits_14_0(mvc_io_wgt_data_bits_14_0),
    .io_wgt_data_bits_14_1(mvc_io_wgt_data_bits_14_1),
    .io_wgt_data_bits_14_2(mvc_io_wgt_data_bits_14_2),
    .io_wgt_data_bits_14_3(mvc_io_wgt_data_bits_14_3),
    .io_wgt_data_bits_14_4(mvc_io_wgt_data_bits_14_4),
    .io_wgt_data_bits_14_5(mvc_io_wgt_data_bits_14_5),
    .io_wgt_data_bits_14_6(mvc_io_wgt_data_bits_14_6),
    .io_wgt_data_bits_14_7(mvc_io_wgt_data_bits_14_7),
    .io_wgt_data_bits_14_8(mvc_io_wgt_data_bits_14_8),
    .io_wgt_data_bits_14_9(mvc_io_wgt_data_bits_14_9),
    .io_wgt_data_bits_14_10(mvc_io_wgt_data_bits_14_10),
    .io_wgt_data_bits_14_11(mvc_io_wgt_data_bits_14_11),
    .io_wgt_data_bits_14_12(mvc_io_wgt_data_bits_14_12),
    .io_wgt_data_bits_14_13(mvc_io_wgt_data_bits_14_13),
    .io_wgt_data_bits_14_14(mvc_io_wgt_data_bits_14_14),
    .io_wgt_data_bits_14_15(mvc_io_wgt_data_bits_14_15),
    .io_wgt_data_bits_15_0(mvc_io_wgt_data_bits_15_0),
    .io_wgt_data_bits_15_1(mvc_io_wgt_data_bits_15_1),
    .io_wgt_data_bits_15_2(mvc_io_wgt_data_bits_15_2),
    .io_wgt_data_bits_15_3(mvc_io_wgt_data_bits_15_3),
    .io_wgt_data_bits_15_4(mvc_io_wgt_data_bits_15_4),
    .io_wgt_data_bits_15_5(mvc_io_wgt_data_bits_15_5),
    .io_wgt_data_bits_15_6(mvc_io_wgt_data_bits_15_6),
    .io_wgt_data_bits_15_7(mvc_io_wgt_data_bits_15_7),
    .io_wgt_data_bits_15_8(mvc_io_wgt_data_bits_15_8),
    .io_wgt_data_bits_15_9(mvc_io_wgt_data_bits_15_9),
    .io_wgt_data_bits_15_10(mvc_io_wgt_data_bits_15_10),
    .io_wgt_data_bits_15_11(mvc_io_wgt_data_bits_15_11),
    .io_wgt_data_bits_15_12(mvc_io_wgt_data_bits_15_12),
    .io_wgt_data_bits_15_13(mvc_io_wgt_data_bits_15_13),
    .io_wgt_data_bits_15_14(mvc_io_wgt_data_bits_15_14),
    .io_wgt_data_bits_15_15(mvc_io_wgt_data_bits_15_15),
    .io_acc_i_data_valid(mvc_io_acc_i_data_valid),
    .io_acc_i_data_bits_0_0(mvc_io_acc_i_data_bits_0_0),
    .io_acc_i_data_bits_0_1(mvc_io_acc_i_data_bits_0_1),
    .io_acc_i_data_bits_0_2(mvc_io_acc_i_data_bits_0_2),
    .io_acc_i_data_bits_0_3(mvc_io_acc_i_data_bits_0_3),
    .io_acc_i_data_bits_0_4(mvc_io_acc_i_data_bits_0_4),
    .io_acc_i_data_bits_0_5(mvc_io_acc_i_data_bits_0_5),
    .io_acc_i_data_bits_0_6(mvc_io_acc_i_data_bits_0_6),
    .io_acc_i_data_bits_0_7(mvc_io_acc_i_data_bits_0_7),
    .io_acc_i_data_bits_0_8(mvc_io_acc_i_data_bits_0_8),
    .io_acc_i_data_bits_0_9(mvc_io_acc_i_data_bits_0_9),
    .io_acc_i_data_bits_0_10(mvc_io_acc_i_data_bits_0_10),
    .io_acc_i_data_bits_0_11(mvc_io_acc_i_data_bits_0_11),
    .io_acc_i_data_bits_0_12(mvc_io_acc_i_data_bits_0_12),
    .io_acc_i_data_bits_0_13(mvc_io_acc_i_data_bits_0_13),
    .io_acc_i_data_bits_0_14(mvc_io_acc_i_data_bits_0_14),
    .io_acc_i_data_bits_0_15(mvc_io_acc_i_data_bits_0_15),
    .io_acc_o_data_valid(mvc_io_acc_o_data_valid),
    .io_acc_o_data_bits_0_0(mvc_io_acc_o_data_bits_0_0),
    .io_acc_o_data_bits_0_1(mvc_io_acc_o_data_bits_0_1),
    .io_acc_o_data_bits_0_2(mvc_io_acc_o_data_bits_0_2),
    .io_acc_o_data_bits_0_3(mvc_io_acc_o_data_bits_0_3),
    .io_acc_o_data_bits_0_4(mvc_io_acc_o_data_bits_0_4),
    .io_acc_o_data_bits_0_5(mvc_io_acc_o_data_bits_0_5),
    .io_acc_o_data_bits_0_6(mvc_io_acc_o_data_bits_0_6),
    .io_acc_o_data_bits_0_7(mvc_io_acc_o_data_bits_0_7),
    .io_acc_o_data_bits_0_8(mvc_io_acc_o_data_bits_0_8),
    .io_acc_o_data_bits_0_9(mvc_io_acc_o_data_bits_0_9),
    .io_acc_o_data_bits_0_10(mvc_io_acc_o_data_bits_0_10),
    .io_acc_o_data_bits_0_11(mvc_io_acc_o_data_bits_0_11),
    .io_acc_o_data_bits_0_12(mvc_io_acc_o_data_bits_0_12),
    .io_acc_o_data_bits_0_13(mvc_io_acc_o_data_bits_0_13),
    .io_acc_o_data_bits_0_14(mvc_io_acc_o_data_bits_0_14),
    .io_acc_o_data_bits_0_15(mvc_io_acc_o_data_bits_0_15),
    .io_out_data_valid(mvc_io_out_data_valid),
    .io_out_data_bits_0_0(mvc_io_out_data_bits_0_0),
    .io_out_data_bits_0_1(mvc_io_out_data_bits_0_1),
    .io_out_data_bits_0_2(mvc_io_out_data_bits_0_2),
    .io_out_data_bits_0_3(mvc_io_out_data_bits_0_3),
    .io_out_data_bits_0_4(mvc_io_out_data_bits_0_4),
    .io_out_data_bits_0_5(mvc_io_out_data_bits_0_5),
    .io_out_data_bits_0_6(mvc_io_out_data_bits_0_6),
    .io_out_data_bits_0_7(mvc_io_out_data_bits_0_7),
    .io_out_data_bits_0_8(mvc_io_out_data_bits_0_8),
    .io_out_data_bits_0_9(mvc_io_out_data_bits_0_9),
    .io_out_data_bits_0_10(mvc_io_out_data_bits_0_10),
    .io_out_data_bits_0_11(mvc_io_out_data_bits_0_11),
    .io_out_data_bits_0_12(mvc_io_out_data_bits_0_12),
    .io_out_data_bits_0_13(mvc_io_out_data_bits_0_13),
    .io_out_data_bits_0_14(mvc_io_out_data_bits_0_14),
    .io_out_data_bits_0_15(mvc_io_out_data_bits_0_15)
  );
  Pipe_16 wrpipe ( // @[TensorGemm.scala 218:22:@20203.4]
    .clock(wrpipe_clock),
    .reset(wrpipe_reset),
    .io_enq_valid(wrpipe_io_enq_valid),
    .io_enq_bits(wrpipe_io_enq_bits),
    .io_deq_valid(wrpipe_io_deq_valid),
    .io_deq_bits(wrpipe_io_deq_bits)
  );
  assign dec_reset = io_inst[7]; // @[TensorGemm.scala 200:29:@20166.4]
  assign dec_uop_begin = io_inst[20:8]; // @[TensorGemm.scala 200:29:@20168.4]
  assign dec_uop_end = io_inst[34:21]; // @[TensorGemm.scala 200:29:@20170.4]
  assign dec_lp_0 = io_inst[48:35]; // @[TensorGemm.scala 200:29:@20172.4]
  assign dec_lp_1 = io_inst[62:49]; // @[TensorGemm.scala 200:29:@20174.4]
  assign dec_acc_0 = io_inst[74:64]; // @[TensorGemm.scala 200:29:@20178.4]
  assign dec_acc_1 = io_inst[85:75]; // @[TensorGemm.scala 200:29:@20180.4]
  assign dec_inp_0 = io_inst[96:86]; // @[TensorGemm.scala 200:29:@20182.4]
  assign dec_inp_1 = io_inst[107:97]; // @[TensorGemm.scala 200:29:@20184.4]
  assign dec_wgt_0 = io_inst[117:108]; // @[TensorGemm.scala 200:29:@20186.4]
  assign dec_wgt_1 = io_inst[127:118]; // @[TensorGemm.scala 200:29:@20188.4]
  assign _T_7688 = inflight == 5'h0; // @[TensorGemm.scala 219:23:@20206.4]
  assign _T_7689 = state == 3'h4; // @[TensorGemm.scala 220:13:@20207.4]
  assign _T_7691 = dec_lp_0 - 14'h1; // @[TensorGemm.scala 221:26:@20208.4]
  assign _T_7692 = $unsigned(_T_7691); // @[TensorGemm.scala 221:26:@20209.4]
  assign _T_7693 = _T_7692[13:0]; // @[TensorGemm.scala 221:26:@20210.4]
  assign _T_7694 = cnt_o == _T_7693; // @[TensorGemm.scala 221:13:@20211.4]
  assign _T_7695 = _T_7689 & _T_7694; // @[TensorGemm.scala 220:22:@20212.4]
  assign _T_7697 = dec_lp_1 - 14'h1; // @[TensorGemm.scala 222:26:@20213.4]
  assign _T_7698 = $unsigned(_T_7697); // @[TensorGemm.scala 222:26:@20214.4]
  assign _T_7699 = _T_7698[13:0]; // @[TensorGemm.scala 222:26:@20215.4]
  assign _T_7700 = cnt_i == _T_7699; // @[TensorGemm.scala 222:13:@20216.4]
  assign _T_7701 = _T_7695 & _T_7700; // @[TensorGemm.scala 221:32:@20217.4]
  assign _T_7703 = dec_uop_end - 14'h1; // @[TensorGemm.scala 223:27:@20218.4]
  assign _T_7704 = $unsigned(_T_7703); // @[TensorGemm.scala 223:27:@20219.4]
  assign _T_7705 = _T_7704[13:0]; // @[TensorGemm.scala 223:27:@20220.4]
  assign _T_7706 = uop_idx == _T_7705; // @[TensorGemm.scala 223:15:@20221.4]
  assign _T_7707 = _T_7701 & _T_7706; // @[TensorGemm.scala 222:32:@20222.4]
  assign _T_7710 = _T_7707 & _T_7688; // @[TensorGemm.scala 223:33:@20224.4]
  assign _T_7711 = state == 3'h5; // @[TensorGemm.scala 225:13:@20225.4]
  assign _T_7712 = _T_7710 | _T_7711; // @[TensorGemm.scala 224:25:@20226.4]
  assign _T_7713 = 3'h0 == state; // @[Conditional.scala 37:30:@20228.4]
  assign _GEN_0 = io_start ? 3'h1 : state; // @[TensorGemm.scala 229:22:@20230.6]
  assign _T_7714 = 3'h1 == state; // @[Conditional.scala 37:30:@20235.6]
  assign _T_7715 = 3'h2 == state; // @[Conditional.scala 37:30:@20240.8]
  assign _T_7716 = 3'h3 == state; // @[Conditional.scala 37:30:@20245.10]
  assign _T_7717 = 3'h4 == state; // @[Conditional.scala 37:30:@20250.12]
  assign _T_7728 = _T_7694 & _T_7700; // @[TensorGemm.scala 244:36:@20260.14]
  assign _T_7734 = _T_7728 & _T_7706; // @[TensorGemm.scala 245:38:@20265.14]
  assign _T_7736 = inflight != 5'h0; // @[TensorGemm.scala 247:23:@20267.16]
  assign _GEN_1 = _T_7736 ? 3'h5 : 3'h0; // @[TensorGemm.scala 247:32:@20268.16]
  assign _GEN_2 = _T_7734 ? _GEN_1 : 3'h1; // @[TensorGemm.scala 246:40:@20266.14]
  assign _T_7737 = 3'h5 == state; // @[Conditional.scala 37:30:@20280.14]
  assign _GEN_3 = _T_7688 ? 3'h0 : state; // @[TensorGemm.scala 257:30:@20283.16]
  assign _GEN_4 = _T_7737 ? _GEN_3 : state; // @[Conditional.scala 39:67:@20281.14]
  assign _GEN_5 = _T_7717 ? _GEN_2 : _GEN_4; // @[Conditional.scala 39:67:@20251.12]
  assign _GEN_6 = _T_7716 ? 3'h4 : _GEN_5; // @[Conditional.scala 39:67:@20246.10]
  assign _GEN_7 = _T_7715 ? 3'h3 : _GEN_6; // @[Conditional.scala 39:67:@20241.8]
  assign _GEN_8 = _T_7714 ? 3'h2 : _GEN_7; // @[Conditional.scala 39:67:@20236.6]
  assign _GEN_9 = _T_7713 ? _GEN_0 : _GEN_8; // @[Conditional.scala 40:58:@20229.4]
  assign _T_7740 = state == 3'h0; // @[TensorGemm.scala 263:14:@20287.4]
  assign _T_7743 = dec_reset == 1'h0; // @[TensorGemm.scala 265:14:@20292.6]
  assign _T_7744 = state == 3'h3; // @[TensorGemm.scala 266:17:@20294.8]
  assign _T_7745 = _T_7744 & mvc_io_acc_o_data_valid; // @[TensorGemm.scala 266:34:@20295.8]
  assign _T_7748 = inflight + 5'h1; // @[TensorGemm.scala 269:28:@20302.12]
  assign _T_7749 = inflight + 5'h1; // @[TensorGemm.scala 269:28:@20303.12]
  assign _T_7751 = inflight - 5'h1; // @[TensorGemm.scala 271:28:@20308.14]
  assign _T_7752 = $unsigned(_T_7751); // @[TensorGemm.scala 271:28:@20309.14]
  assign _T_7753 = _T_7752[4:0]; // @[TensorGemm.scala 271:28:@20310.14]
  assign _GEN_10 = mvc_io_acc_o_data_valid ? _T_7753 : inflight; // @[TensorGemm.scala 270:41:@20307.12]
  assign _GEN_11 = _T_7744 ? _T_7749 : _GEN_10; // @[TensorGemm.scala 268:39:@20301.10]
  assign _GEN_12 = _T_7745 ? inflight : _GEN_11; // @[TensorGemm.scala 266:62:@20296.8]
  assign _GEN_13 = _T_7743 ? _GEN_12 : inflight; // @[TensorGemm.scala 265:26:@20293.6]
  assign _T_7761 = _T_7689 & _T_7706; // @[TensorGemm.scala 277:23:@20320.4]
  assign _T_7762 = _T_7740 | _T_7761; // @[TensorGemm.scala 276:21:@20321.4]
  assign _GEN_40 = {{1'd0}, dec_uop_begin}; // @[TensorGemm.scala 280:46:@20327.6]
  assign _T_7764 = _GEN_40 != dec_uop_end; // @[TensorGemm.scala 280:46:@20327.6]
  assign _T_7765 = _T_7689 & _T_7764; // @[TensorGemm.scala 280:29:@20328.6]
  assign _T_7767 = uop_idx + 14'h1; // @[TensorGemm.scala 281:24:@20330.8]
  assign _T_7768 = uop_idx + 14'h1; // @[TensorGemm.scala 281:24:@20331.8]
  assign _GEN_15 = _T_7765 ? _T_7768 : uop_idx; // @[TensorGemm.scala 280:59:@20329.6]
  assign _T_7786 = _T_7761 & _T_7700; // @[TensorGemm.scala 291:33:@20352.6]
  assign _T_7788 = cnt_o + 14'h1; // @[TensorGemm.scala 293:20:@20354.8]
  assign _T_7789 = cnt_o + 14'h1; // @[TensorGemm.scala 293:20:@20355.8]
  assign _GEN_41 = {{3'd0}, dec_acc_0}; // @[TensorGemm.scala 294:20:@20357.8]
  assign _T_7790 = acc_o + _GEN_41; // @[TensorGemm.scala 294:20:@20357.8]
  assign _T_7791 = acc_o + _GEN_41; // @[TensorGemm.scala 294:20:@20358.8]
  assign _GEN_42 = {{3'd0}, dec_inp_0}; // @[TensorGemm.scala 295:20:@20360.8]
  assign _T_7792 = inp_o + _GEN_42; // @[TensorGemm.scala 295:20:@20360.8]
  assign _T_7793 = inp_o + _GEN_42; // @[TensorGemm.scala 295:20:@20361.8]
  assign _GEN_43 = {{4'd0}, dec_wgt_0}; // @[TensorGemm.scala 296:20:@20363.8]
  assign _T_7794 = wgt_o + _GEN_43; // @[TensorGemm.scala 296:20:@20363.8]
  assign _T_7795 = wgt_o + _GEN_43; // @[TensorGemm.scala 296:20:@20364.8]
  assign _GEN_17 = _T_7786 ? _T_7789 : cnt_o; // @[TensorGemm.scala 292:33:@20353.6]
  assign _GEN_18 = _T_7786 ? _T_7791 : acc_o; // @[TensorGemm.scala 292:33:@20353.6]
  assign _GEN_19 = _T_7786 ? _T_7793 : inp_o; // @[TensorGemm.scala 292:33:@20353.6]
  assign _GEN_20 = _T_7786 ? _T_7795 : wgt_o; // @[TensorGemm.scala 292:33:@20353.6]
  assign _T_7801 = state == 3'h1; // @[TensorGemm.scala 304:20:@20375.6]
  assign _T_7802 = cnt_i == dec_lp_1; // @[TensorGemm.scala 304:42:@20376.6]
  assign _T_7803 = _T_7801 & _T_7802; // @[TensorGemm.scala 304:33:@20377.6]
  assign _T_7813 = cnt_i + 14'h1; // @[TensorGemm.scala 310:20:@20392.10]
  assign _T_7814 = cnt_i + 14'h1; // @[TensorGemm.scala 310:20:@20393.10]
  assign _GEN_44 = {{3'd0}, dec_acc_1}; // @[TensorGemm.scala 311:20:@20395.10]
  assign _T_7815 = acc_i + _GEN_44; // @[TensorGemm.scala 311:20:@20395.10]
  assign _T_7816 = acc_i + _GEN_44; // @[TensorGemm.scala 311:20:@20396.10]
  assign _GEN_45 = {{3'd0}, dec_inp_1}; // @[TensorGemm.scala 312:20:@20398.10]
  assign _T_7817 = inp_i + _GEN_45; // @[TensorGemm.scala 312:20:@20398.10]
  assign _T_7818 = inp_i + _GEN_45; // @[TensorGemm.scala 312:20:@20399.10]
  assign _GEN_46 = {{4'd0}, dec_wgt_1}; // @[TensorGemm.scala 313:20:@20401.10]
  assign _T_7819 = wgt_i + _GEN_46; // @[TensorGemm.scala 313:20:@20401.10]
  assign _T_7820 = wgt_i + _GEN_46; // @[TensorGemm.scala 313:20:@20402.10]
  assign _GEN_25 = _T_7761 ? _T_7814 : cnt_i; // @[TensorGemm.scala 309:59:@20391.8]
  assign _GEN_26 = _T_7761 ? _T_7816 : acc_i; // @[TensorGemm.scala 309:59:@20391.8]
  assign _GEN_27 = _T_7761 ? _T_7818 : inp_i; // @[TensorGemm.scala 309:59:@20391.8]
  assign _GEN_28 = _T_7761 ? _T_7820 : wgt_i; // @[TensorGemm.scala 309:59:@20391.8]
  assign _GEN_29 = _T_7803 ? 14'h0 : _GEN_25; // @[TensorGemm.scala 304:56:@20378.6]
  assign _GEN_30 = _T_7803 ? acc_o : _GEN_26; // @[TensorGemm.scala 304:56:@20378.6]
  assign _GEN_31 = _T_7803 ? inp_o : _GEN_27; // @[TensorGemm.scala 304:56:@20378.6]
  assign _GEN_32 = _T_7803 ? wgt_o : _GEN_28; // @[TensorGemm.scala 304:56:@20378.6]
  assign _T_7821 = state == 3'h2; // @[TensorGemm.scala 316:14:@20405.4]
  assign _T_7822 = _T_7821 & io_uop_data_valid; // @[TensorGemm.scala 316:30:@20406.4]
  assign _GEN_47 = {{3'd0}, io_uop_data_bits_u0}; // @[TensorGemm.scala 317:36:@20408.6]
  assign _T_7823 = _GEN_47 + acc_i; // @[TensorGemm.scala 317:36:@20408.6]
  assign _T_7824 = _GEN_47 + acc_i; // @[TensorGemm.scala 317:36:@20409.6]
  assign _GEN_48 = {{3'd0}, io_uop_data_bits_u1}; // @[TensorGemm.scala 318:36:@20411.6]
  assign _T_7825 = _GEN_48 + inp_i; // @[TensorGemm.scala 318:36:@20411.6]
  assign _T_7826 = _GEN_48 + inp_i; // @[TensorGemm.scala 318:36:@20412.6]
  assign _GEN_49 = {{4'd0}, io_uop_data_bits_u2}; // @[TensorGemm.scala 319:36:@20414.6]
  assign _T_7827 = _GEN_49 + wgt_i; // @[TensorGemm.scala 319:36:@20414.6]
  assign _T_7828 = _GEN_49 + wgt_i; // @[TensorGemm.scala 319:36:@20415.6]
  assign _T_7830 = ~ dec_reset; // @[TensorGemm.scala 322:43:@20419.4]
  assign _T_8115 = dec_reset ? 1'h1 : wrpipe_io_deq_valid; // @[TensorGemm.scala 351:8:@21005.4]
  assign _T_8117 = dec_reset ? uop_acc : wrpipe_io_deq_bits; // @[TensorGemm.scala 352:28:@21008.4]
  assign io_done = _T_7688 & _T_7712; // @[TensorGemm.scala 361:11:@21047.4]
  assign io_uop_idx_valid = state == 3'h1; // @[TensorGemm.scala 326:20:@20424.4]
  assign io_uop_idx_bits = uop_idx[10:0]; // @[TensorGemm.scala 327:19:@20425.4]
  assign io_inp_rd_idx_valid = state == 3'h3; // @[TensorGemm.scala 330:23:@20427.4]
  assign io_inp_rd_idx_bits = uop_inp[10:0]; // @[TensorGemm.scala 331:22:@20428.4]
  assign io_wgt_rd_idx_valid = state == 3'h3; // @[TensorGemm.scala 335:23:@20448.4]
  assign io_wgt_rd_idx_bits = uop_wgt[9:0]; // @[TensorGemm.scala 336:22:@20449.4]
  assign io_acc_rd_idx_valid = state == 3'h3; // @[TensorGemm.scala 340:23:@20709.4]
  assign io_acc_rd_idx_bits = uop_acc[10:0]; // @[TensorGemm.scala 341:22:@20710.4]
  assign io_acc_wr_valid = mvc_io_acc_o_data_valid & _T_8115; // @[TensorGemm.scala 350:19:@21007.4]
  assign io_acc_wr_bits_idx = _T_8117[10:0]; // @[TensorGemm.scala 352:22:@21009.4]
  assign io_acc_wr_bits_data_0_0 = mvc_io_acc_o_data_bits_0_0; // @[TensorGemm.scala 353:23:@21010.4]
  assign io_acc_wr_bits_data_0_1 = mvc_io_acc_o_data_bits_0_1; // @[TensorGemm.scala 353:23:@21011.4]
  assign io_acc_wr_bits_data_0_2 = mvc_io_acc_o_data_bits_0_2; // @[TensorGemm.scala 353:23:@21012.4]
  assign io_acc_wr_bits_data_0_3 = mvc_io_acc_o_data_bits_0_3; // @[TensorGemm.scala 353:23:@21013.4]
  assign io_acc_wr_bits_data_0_4 = mvc_io_acc_o_data_bits_0_4; // @[TensorGemm.scala 353:23:@21014.4]
  assign io_acc_wr_bits_data_0_5 = mvc_io_acc_o_data_bits_0_5; // @[TensorGemm.scala 353:23:@21015.4]
  assign io_acc_wr_bits_data_0_6 = mvc_io_acc_o_data_bits_0_6; // @[TensorGemm.scala 353:23:@21016.4]
  assign io_acc_wr_bits_data_0_7 = mvc_io_acc_o_data_bits_0_7; // @[TensorGemm.scala 353:23:@21017.4]
  assign io_acc_wr_bits_data_0_8 = mvc_io_acc_o_data_bits_0_8; // @[TensorGemm.scala 353:23:@21018.4]
  assign io_acc_wr_bits_data_0_9 = mvc_io_acc_o_data_bits_0_9; // @[TensorGemm.scala 353:23:@21019.4]
  assign io_acc_wr_bits_data_0_10 = mvc_io_acc_o_data_bits_0_10; // @[TensorGemm.scala 353:23:@21020.4]
  assign io_acc_wr_bits_data_0_11 = mvc_io_acc_o_data_bits_0_11; // @[TensorGemm.scala 353:23:@21021.4]
  assign io_acc_wr_bits_data_0_12 = mvc_io_acc_o_data_bits_0_12; // @[TensorGemm.scala 353:23:@21022.4]
  assign io_acc_wr_bits_data_0_13 = mvc_io_acc_o_data_bits_0_13; // @[TensorGemm.scala 353:23:@21023.4]
  assign io_acc_wr_bits_data_0_14 = mvc_io_acc_o_data_bits_0_14; // @[TensorGemm.scala 353:23:@21024.4]
  assign io_acc_wr_bits_data_0_15 = mvc_io_acc_o_data_bits_0_15; // @[TensorGemm.scala 353:23:@21025.4]
  assign io_out_wr_valid = mvc_io_out_data_valid & wrpipe_io_deq_valid; // @[TensorGemm.scala 356:19:@21027.4]
  assign io_out_wr_bits_idx = wrpipe_io_deq_bits[10:0]; // @[TensorGemm.scala 357:22:@21028.4]
  assign io_out_wr_bits_data_0_0 = mvc_io_out_data_bits_0_0; // @[TensorGemm.scala 358:23:@21029.4]
  assign io_out_wr_bits_data_0_1 = mvc_io_out_data_bits_0_1; // @[TensorGemm.scala 358:23:@21030.4]
  assign io_out_wr_bits_data_0_2 = mvc_io_out_data_bits_0_2; // @[TensorGemm.scala 358:23:@21031.4]
  assign io_out_wr_bits_data_0_3 = mvc_io_out_data_bits_0_3; // @[TensorGemm.scala 358:23:@21032.4]
  assign io_out_wr_bits_data_0_4 = mvc_io_out_data_bits_0_4; // @[TensorGemm.scala 358:23:@21033.4]
  assign io_out_wr_bits_data_0_5 = mvc_io_out_data_bits_0_5; // @[TensorGemm.scala 358:23:@21034.4]
  assign io_out_wr_bits_data_0_6 = mvc_io_out_data_bits_0_6; // @[TensorGemm.scala 358:23:@21035.4]
  assign io_out_wr_bits_data_0_7 = mvc_io_out_data_bits_0_7; // @[TensorGemm.scala 358:23:@21036.4]
  assign io_out_wr_bits_data_0_8 = mvc_io_out_data_bits_0_8; // @[TensorGemm.scala 358:23:@21037.4]
  assign io_out_wr_bits_data_0_9 = mvc_io_out_data_bits_0_9; // @[TensorGemm.scala 358:23:@21038.4]
  assign io_out_wr_bits_data_0_10 = mvc_io_out_data_bits_0_10; // @[TensorGemm.scala 358:23:@21039.4]
  assign io_out_wr_bits_data_0_11 = mvc_io_out_data_bits_0_11; // @[TensorGemm.scala 358:23:@21040.4]
  assign io_out_wr_bits_data_0_12 = mvc_io_out_data_bits_0_12; // @[TensorGemm.scala 358:23:@21041.4]
  assign io_out_wr_bits_data_0_13 = mvc_io_out_data_bits_0_13; // @[TensorGemm.scala 358:23:@21042.4]
  assign io_out_wr_bits_data_0_14 = mvc_io_out_data_bits_0_14; // @[TensorGemm.scala 358:23:@21043.4]
  assign io_out_wr_bits_data_0_15 = mvc_io_out_data_bits_0_15; // @[TensorGemm.scala 358:23:@21044.4]
  assign mvc_clock = clock; // @[:@20151.4]
  assign mvc_reset = reset; // @[:@20152.4]
  assign mvc_io_reset = dec_reset & _T_7689; // @[TensorGemm.scala 344:16:@20713.4]
  assign mvc_io_inp_data_valid = io_inp_rd_data_valid; // @[TensorGemm.scala 345:19:@20730.4]
  assign mvc_io_inp_data_bits_0_0 = io_inp_rd_data_bits_0_0; // @[TensorGemm.scala 345:19:@20714.4]
  assign mvc_io_inp_data_bits_0_1 = io_inp_rd_data_bits_0_1; // @[TensorGemm.scala 345:19:@20715.4]
  assign mvc_io_inp_data_bits_0_2 = io_inp_rd_data_bits_0_2; // @[TensorGemm.scala 345:19:@20716.4]
  assign mvc_io_inp_data_bits_0_3 = io_inp_rd_data_bits_0_3; // @[TensorGemm.scala 345:19:@20717.4]
  assign mvc_io_inp_data_bits_0_4 = io_inp_rd_data_bits_0_4; // @[TensorGemm.scala 345:19:@20718.4]
  assign mvc_io_inp_data_bits_0_5 = io_inp_rd_data_bits_0_5; // @[TensorGemm.scala 345:19:@20719.4]
  assign mvc_io_inp_data_bits_0_6 = io_inp_rd_data_bits_0_6; // @[TensorGemm.scala 345:19:@20720.4]
  assign mvc_io_inp_data_bits_0_7 = io_inp_rd_data_bits_0_7; // @[TensorGemm.scala 345:19:@20721.4]
  assign mvc_io_inp_data_bits_0_8 = io_inp_rd_data_bits_0_8; // @[TensorGemm.scala 345:19:@20722.4]
  assign mvc_io_inp_data_bits_0_9 = io_inp_rd_data_bits_0_9; // @[TensorGemm.scala 345:19:@20723.4]
  assign mvc_io_inp_data_bits_0_10 = io_inp_rd_data_bits_0_10; // @[TensorGemm.scala 345:19:@20724.4]
  assign mvc_io_inp_data_bits_0_11 = io_inp_rd_data_bits_0_11; // @[TensorGemm.scala 345:19:@20725.4]
  assign mvc_io_inp_data_bits_0_12 = io_inp_rd_data_bits_0_12; // @[TensorGemm.scala 345:19:@20726.4]
  assign mvc_io_inp_data_bits_0_13 = io_inp_rd_data_bits_0_13; // @[TensorGemm.scala 345:19:@20727.4]
  assign mvc_io_inp_data_bits_0_14 = io_inp_rd_data_bits_0_14; // @[TensorGemm.scala 345:19:@20728.4]
  assign mvc_io_inp_data_bits_0_15 = io_inp_rd_data_bits_0_15; // @[TensorGemm.scala 345:19:@20729.4]
  assign mvc_io_wgt_data_valid = io_wgt_rd_data_valid; // @[TensorGemm.scala 346:19:@20987.4]
  assign mvc_io_wgt_data_bits_0_0 = io_wgt_rd_data_bits_0_0; // @[TensorGemm.scala 346:19:@20731.4]
  assign mvc_io_wgt_data_bits_0_1 = io_wgt_rd_data_bits_0_1; // @[TensorGemm.scala 346:19:@20732.4]
  assign mvc_io_wgt_data_bits_0_2 = io_wgt_rd_data_bits_0_2; // @[TensorGemm.scala 346:19:@20733.4]
  assign mvc_io_wgt_data_bits_0_3 = io_wgt_rd_data_bits_0_3; // @[TensorGemm.scala 346:19:@20734.4]
  assign mvc_io_wgt_data_bits_0_4 = io_wgt_rd_data_bits_0_4; // @[TensorGemm.scala 346:19:@20735.4]
  assign mvc_io_wgt_data_bits_0_5 = io_wgt_rd_data_bits_0_5; // @[TensorGemm.scala 346:19:@20736.4]
  assign mvc_io_wgt_data_bits_0_6 = io_wgt_rd_data_bits_0_6; // @[TensorGemm.scala 346:19:@20737.4]
  assign mvc_io_wgt_data_bits_0_7 = io_wgt_rd_data_bits_0_7; // @[TensorGemm.scala 346:19:@20738.4]
  assign mvc_io_wgt_data_bits_0_8 = io_wgt_rd_data_bits_0_8; // @[TensorGemm.scala 346:19:@20739.4]
  assign mvc_io_wgt_data_bits_0_9 = io_wgt_rd_data_bits_0_9; // @[TensorGemm.scala 346:19:@20740.4]
  assign mvc_io_wgt_data_bits_0_10 = io_wgt_rd_data_bits_0_10; // @[TensorGemm.scala 346:19:@20741.4]
  assign mvc_io_wgt_data_bits_0_11 = io_wgt_rd_data_bits_0_11; // @[TensorGemm.scala 346:19:@20742.4]
  assign mvc_io_wgt_data_bits_0_12 = io_wgt_rd_data_bits_0_12; // @[TensorGemm.scala 346:19:@20743.4]
  assign mvc_io_wgt_data_bits_0_13 = io_wgt_rd_data_bits_0_13; // @[TensorGemm.scala 346:19:@20744.4]
  assign mvc_io_wgt_data_bits_0_14 = io_wgt_rd_data_bits_0_14; // @[TensorGemm.scala 346:19:@20745.4]
  assign mvc_io_wgt_data_bits_0_15 = io_wgt_rd_data_bits_0_15; // @[TensorGemm.scala 346:19:@20746.4]
  assign mvc_io_wgt_data_bits_1_0 = io_wgt_rd_data_bits_1_0; // @[TensorGemm.scala 346:19:@20747.4]
  assign mvc_io_wgt_data_bits_1_1 = io_wgt_rd_data_bits_1_1; // @[TensorGemm.scala 346:19:@20748.4]
  assign mvc_io_wgt_data_bits_1_2 = io_wgt_rd_data_bits_1_2; // @[TensorGemm.scala 346:19:@20749.4]
  assign mvc_io_wgt_data_bits_1_3 = io_wgt_rd_data_bits_1_3; // @[TensorGemm.scala 346:19:@20750.4]
  assign mvc_io_wgt_data_bits_1_4 = io_wgt_rd_data_bits_1_4; // @[TensorGemm.scala 346:19:@20751.4]
  assign mvc_io_wgt_data_bits_1_5 = io_wgt_rd_data_bits_1_5; // @[TensorGemm.scala 346:19:@20752.4]
  assign mvc_io_wgt_data_bits_1_6 = io_wgt_rd_data_bits_1_6; // @[TensorGemm.scala 346:19:@20753.4]
  assign mvc_io_wgt_data_bits_1_7 = io_wgt_rd_data_bits_1_7; // @[TensorGemm.scala 346:19:@20754.4]
  assign mvc_io_wgt_data_bits_1_8 = io_wgt_rd_data_bits_1_8; // @[TensorGemm.scala 346:19:@20755.4]
  assign mvc_io_wgt_data_bits_1_9 = io_wgt_rd_data_bits_1_9; // @[TensorGemm.scala 346:19:@20756.4]
  assign mvc_io_wgt_data_bits_1_10 = io_wgt_rd_data_bits_1_10; // @[TensorGemm.scala 346:19:@20757.4]
  assign mvc_io_wgt_data_bits_1_11 = io_wgt_rd_data_bits_1_11; // @[TensorGemm.scala 346:19:@20758.4]
  assign mvc_io_wgt_data_bits_1_12 = io_wgt_rd_data_bits_1_12; // @[TensorGemm.scala 346:19:@20759.4]
  assign mvc_io_wgt_data_bits_1_13 = io_wgt_rd_data_bits_1_13; // @[TensorGemm.scala 346:19:@20760.4]
  assign mvc_io_wgt_data_bits_1_14 = io_wgt_rd_data_bits_1_14; // @[TensorGemm.scala 346:19:@20761.4]
  assign mvc_io_wgt_data_bits_1_15 = io_wgt_rd_data_bits_1_15; // @[TensorGemm.scala 346:19:@20762.4]
  assign mvc_io_wgt_data_bits_2_0 = io_wgt_rd_data_bits_2_0; // @[TensorGemm.scala 346:19:@20763.4]
  assign mvc_io_wgt_data_bits_2_1 = io_wgt_rd_data_bits_2_1; // @[TensorGemm.scala 346:19:@20764.4]
  assign mvc_io_wgt_data_bits_2_2 = io_wgt_rd_data_bits_2_2; // @[TensorGemm.scala 346:19:@20765.4]
  assign mvc_io_wgt_data_bits_2_3 = io_wgt_rd_data_bits_2_3; // @[TensorGemm.scala 346:19:@20766.4]
  assign mvc_io_wgt_data_bits_2_4 = io_wgt_rd_data_bits_2_4; // @[TensorGemm.scala 346:19:@20767.4]
  assign mvc_io_wgt_data_bits_2_5 = io_wgt_rd_data_bits_2_5; // @[TensorGemm.scala 346:19:@20768.4]
  assign mvc_io_wgt_data_bits_2_6 = io_wgt_rd_data_bits_2_6; // @[TensorGemm.scala 346:19:@20769.4]
  assign mvc_io_wgt_data_bits_2_7 = io_wgt_rd_data_bits_2_7; // @[TensorGemm.scala 346:19:@20770.4]
  assign mvc_io_wgt_data_bits_2_8 = io_wgt_rd_data_bits_2_8; // @[TensorGemm.scala 346:19:@20771.4]
  assign mvc_io_wgt_data_bits_2_9 = io_wgt_rd_data_bits_2_9; // @[TensorGemm.scala 346:19:@20772.4]
  assign mvc_io_wgt_data_bits_2_10 = io_wgt_rd_data_bits_2_10; // @[TensorGemm.scala 346:19:@20773.4]
  assign mvc_io_wgt_data_bits_2_11 = io_wgt_rd_data_bits_2_11; // @[TensorGemm.scala 346:19:@20774.4]
  assign mvc_io_wgt_data_bits_2_12 = io_wgt_rd_data_bits_2_12; // @[TensorGemm.scala 346:19:@20775.4]
  assign mvc_io_wgt_data_bits_2_13 = io_wgt_rd_data_bits_2_13; // @[TensorGemm.scala 346:19:@20776.4]
  assign mvc_io_wgt_data_bits_2_14 = io_wgt_rd_data_bits_2_14; // @[TensorGemm.scala 346:19:@20777.4]
  assign mvc_io_wgt_data_bits_2_15 = io_wgt_rd_data_bits_2_15; // @[TensorGemm.scala 346:19:@20778.4]
  assign mvc_io_wgt_data_bits_3_0 = io_wgt_rd_data_bits_3_0; // @[TensorGemm.scala 346:19:@20779.4]
  assign mvc_io_wgt_data_bits_3_1 = io_wgt_rd_data_bits_3_1; // @[TensorGemm.scala 346:19:@20780.4]
  assign mvc_io_wgt_data_bits_3_2 = io_wgt_rd_data_bits_3_2; // @[TensorGemm.scala 346:19:@20781.4]
  assign mvc_io_wgt_data_bits_3_3 = io_wgt_rd_data_bits_3_3; // @[TensorGemm.scala 346:19:@20782.4]
  assign mvc_io_wgt_data_bits_3_4 = io_wgt_rd_data_bits_3_4; // @[TensorGemm.scala 346:19:@20783.4]
  assign mvc_io_wgt_data_bits_3_5 = io_wgt_rd_data_bits_3_5; // @[TensorGemm.scala 346:19:@20784.4]
  assign mvc_io_wgt_data_bits_3_6 = io_wgt_rd_data_bits_3_6; // @[TensorGemm.scala 346:19:@20785.4]
  assign mvc_io_wgt_data_bits_3_7 = io_wgt_rd_data_bits_3_7; // @[TensorGemm.scala 346:19:@20786.4]
  assign mvc_io_wgt_data_bits_3_8 = io_wgt_rd_data_bits_3_8; // @[TensorGemm.scala 346:19:@20787.4]
  assign mvc_io_wgt_data_bits_3_9 = io_wgt_rd_data_bits_3_9; // @[TensorGemm.scala 346:19:@20788.4]
  assign mvc_io_wgt_data_bits_3_10 = io_wgt_rd_data_bits_3_10; // @[TensorGemm.scala 346:19:@20789.4]
  assign mvc_io_wgt_data_bits_3_11 = io_wgt_rd_data_bits_3_11; // @[TensorGemm.scala 346:19:@20790.4]
  assign mvc_io_wgt_data_bits_3_12 = io_wgt_rd_data_bits_3_12; // @[TensorGemm.scala 346:19:@20791.4]
  assign mvc_io_wgt_data_bits_3_13 = io_wgt_rd_data_bits_3_13; // @[TensorGemm.scala 346:19:@20792.4]
  assign mvc_io_wgt_data_bits_3_14 = io_wgt_rd_data_bits_3_14; // @[TensorGemm.scala 346:19:@20793.4]
  assign mvc_io_wgt_data_bits_3_15 = io_wgt_rd_data_bits_3_15; // @[TensorGemm.scala 346:19:@20794.4]
  assign mvc_io_wgt_data_bits_4_0 = io_wgt_rd_data_bits_4_0; // @[TensorGemm.scala 346:19:@20795.4]
  assign mvc_io_wgt_data_bits_4_1 = io_wgt_rd_data_bits_4_1; // @[TensorGemm.scala 346:19:@20796.4]
  assign mvc_io_wgt_data_bits_4_2 = io_wgt_rd_data_bits_4_2; // @[TensorGemm.scala 346:19:@20797.4]
  assign mvc_io_wgt_data_bits_4_3 = io_wgt_rd_data_bits_4_3; // @[TensorGemm.scala 346:19:@20798.4]
  assign mvc_io_wgt_data_bits_4_4 = io_wgt_rd_data_bits_4_4; // @[TensorGemm.scala 346:19:@20799.4]
  assign mvc_io_wgt_data_bits_4_5 = io_wgt_rd_data_bits_4_5; // @[TensorGemm.scala 346:19:@20800.4]
  assign mvc_io_wgt_data_bits_4_6 = io_wgt_rd_data_bits_4_6; // @[TensorGemm.scala 346:19:@20801.4]
  assign mvc_io_wgt_data_bits_4_7 = io_wgt_rd_data_bits_4_7; // @[TensorGemm.scala 346:19:@20802.4]
  assign mvc_io_wgt_data_bits_4_8 = io_wgt_rd_data_bits_4_8; // @[TensorGemm.scala 346:19:@20803.4]
  assign mvc_io_wgt_data_bits_4_9 = io_wgt_rd_data_bits_4_9; // @[TensorGemm.scala 346:19:@20804.4]
  assign mvc_io_wgt_data_bits_4_10 = io_wgt_rd_data_bits_4_10; // @[TensorGemm.scala 346:19:@20805.4]
  assign mvc_io_wgt_data_bits_4_11 = io_wgt_rd_data_bits_4_11; // @[TensorGemm.scala 346:19:@20806.4]
  assign mvc_io_wgt_data_bits_4_12 = io_wgt_rd_data_bits_4_12; // @[TensorGemm.scala 346:19:@20807.4]
  assign mvc_io_wgt_data_bits_4_13 = io_wgt_rd_data_bits_4_13; // @[TensorGemm.scala 346:19:@20808.4]
  assign mvc_io_wgt_data_bits_4_14 = io_wgt_rd_data_bits_4_14; // @[TensorGemm.scala 346:19:@20809.4]
  assign mvc_io_wgt_data_bits_4_15 = io_wgt_rd_data_bits_4_15; // @[TensorGemm.scala 346:19:@20810.4]
  assign mvc_io_wgt_data_bits_5_0 = io_wgt_rd_data_bits_5_0; // @[TensorGemm.scala 346:19:@20811.4]
  assign mvc_io_wgt_data_bits_5_1 = io_wgt_rd_data_bits_5_1; // @[TensorGemm.scala 346:19:@20812.4]
  assign mvc_io_wgt_data_bits_5_2 = io_wgt_rd_data_bits_5_2; // @[TensorGemm.scala 346:19:@20813.4]
  assign mvc_io_wgt_data_bits_5_3 = io_wgt_rd_data_bits_5_3; // @[TensorGemm.scala 346:19:@20814.4]
  assign mvc_io_wgt_data_bits_5_4 = io_wgt_rd_data_bits_5_4; // @[TensorGemm.scala 346:19:@20815.4]
  assign mvc_io_wgt_data_bits_5_5 = io_wgt_rd_data_bits_5_5; // @[TensorGemm.scala 346:19:@20816.4]
  assign mvc_io_wgt_data_bits_5_6 = io_wgt_rd_data_bits_5_6; // @[TensorGemm.scala 346:19:@20817.4]
  assign mvc_io_wgt_data_bits_5_7 = io_wgt_rd_data_bits_5_7; // @[TensorGemm.scala 346:19:@20818.4]
  assign mvc_io_wgt_data_bits_5_8 = io_wgt_rd_data_bits_5_8; // @[TensorGemm.scala 346:19:@20819.4]
  assign mvc_io_wgt_data_bits_5_9 = io_wgt_rd_data_bits_5_9; // @[TensorGemm.scala 346:19:@20820.4]
  assign mvc_io_wgt_data_bits_5_10 = io_wgt_rd_data_bits_5_10; // @[TensorGemm.scala 346:19:@20821.4]
  assign mvc_io_wgt_data_bits_5_11 = io_wgt_rd_data_bits_5_11; // @[TensorGemm.scala 346:19:@20822.4]
  assign mvc_io_wgt_data_bits_5_12 = io_wgt_rd_data_bits_5_12; // @[TensorGemm.scala 346:19:@20823.4]
  assign mvc_io_wgt_data_bits_5_13 = io_wgt_rd_data_bits_5_13; // @[TensorGemm.scala 346:19:@20824.4]
  assign mvc_io_wgt_data_bits_5_14 = io_wgt_rd_data_bits_5_14; // @[TensorGemm.scala 346:19:@20825.4]
  assign mvc_io_wgt_data_bits_5_15 = io_wgt_rd_data_bits_5_15; // @[TensorGemm.scala 346:19:@20826.4]
  assign mvc_io_wgt_data_bits_6_0 = io_wgt_rd_data_bits_6_0; // @[TensorGemm.scala 346:19:@20827.4]
  assign mvc_io_wgt_data_bits_6_1 = io_wgt_rd_data_bits_6_1; // @[TensorGemm.scala 346:19:@20828.4]
  assign mvc_io_wgt_data_bits_6_2 = io_wgt_rd_data_bits_6_2; // @[TensorGemm.scala 346:19:@20829.4]
  assign mvc_io_wgt_data_bits_6_3 = io_wgt_rd_data_bits_6_3; // @[TensorGemm.scala 346:19:@20830.4]
  assign mvc_io_wgt_data_bits_6_4 = io_wgt_rd_data_bits_6_4; // @[TensorGemm.scala 346:19:@20831.4]
  assign mvc_io_wgt_data_bits_6_5 = io_wgt_rd_data_bits_6_5; // @[TensorGemm.scala 346:19:@20832.4]
  assign mvc_io_wgt_data_bits_6_6 = io_wgt_rd_data_bits_6_6; // @[TensorGemm.scala 346:19:@20833.4]
  assign mvc_io_wgt_data_bits_6_7 = io_wgt_rd_data_bits_6_7; // @[TensorGemm.scala 346:19:@20834.4]
  assign mvc_io_wgt_data_bits_6_8 = io_wgt_rd_data_bits_6_8; // @[TensorGemm.scala 346:19:@20835.4]
  assign mvc_io_wgt_data_bits_6_9 = io_wgt_rd_data_bits_6_9; // @[TensorGemm.scala 346:19:@20836.4]
  assign mvc_io_wgt_data_bits_6_10 = io_wgt_rd_data_bits_6_10; // @[TensorGemm.scala 346:19:@20837.4]
  assign mvc_io_wgt_data_bits_6_11 = io_wgt_rd_data_bits_6_11; // @[TensorGemm.scala 346:19:@20838.4]
  assign mvc_io_wgt_data_bits_6_12 = io_wgt_rd_data_bits_6_12; // @[TensorGemm.scala 346:19:@20839.4]
  assign mvc_io_wgt_data_bits_6_13 = io_wgt_rd_data_bits_6_13; // @[TensorGemm.scala 346:19:@20840.4]
  assign mvc_io_wgt_data_bits_6_14 = io_wgt_rd_data_bits_6_14; // @[TensorGemm.scala 346:19:@20841.4]
  assign mvc_io_wgt_data_bits_6_15 = io_wgt_rd_data_bits_6_15; // @[TensorGemm.scala 346:19:@20842.4]
  assign mvc_io_wgt_data_bits_7_0 = io_wgt_rd_data_bits_7_0; // @[TensorGemm.scala 346:19:@20843.4]
  assign mvc_io_wgt_data_bits_7_1 = io_wgt_rd_data_bits_7_1; // @[TensorGemm.scala 346:19:@20844.4]
  assign mvc_io_wgt_data_bits_7_2 = io_wgt_rd_data_bits_7_2; // @[TensorGemm.scala 346:19:@20845.4]
  assign mvc_io_wgt_data_bits_7_3 = io_wgt_rd_data_bits_7_3; // @[TensorGemm.scala 346:19:@20846.4]
  assign mvc_io_wgt_data_bits_7_4 = io_wgt_rd_data_bits_7_4; // @[TensorGemm.scala 346:19:@20847.4]
  assign mvc_io_wgt_data_bits_7_5 = io_wgt_rd_data_bits_7_5; // @[TensorGemm.scala 346:19:@20848.4]
  assign mvc_io_wgt_data_bits_7_6 = io_wgt_rd_data_bits_7_6; // @[TensorGemm.scala 346:19:@20849.4]
  assign mvc_io_wgt_data_bits_7_7 = io_wgt_rd_data_bits_7_7; // @[TensorGemm.scala 346:19:@20850.4]
  assign mvc_io_wgt_data_bits_7_8 = io_wgt_rd_data_bits_7_8; // @[TensorGemm.scala 346:19:@20851.4]
  assign mvc_io_wgt_data_bits_7_9 = io_wgt_rd_data_bits_7_9; // @[TensorGemm.scala 346:19:@20852.4]
  assign mvc_io_wgt_data_bits_7_10 = io_wgt_rd_data_bits_7_10; // @[TensorGemm.scala 346:19:@20853.4]
  assign mvc_io_wgt_data_bits_7_11 = io_wgt_rd_data_bits_7_11; // @[TensorGemm.scala 346:19:@20854.4]
  assign mvc_io_wgt_data_bits_7_12 = io_wgt_rd_data_bits_7_12; // @[TensorGemm.scala 346:19:@20855.4]
  assign mvc_io_wgt_data_bits_7_13 = io_wgt_rd_data_bits_7_13; // @[TensorGemm.scala 346:19:@20856.4]
  assign mvc_io_wgt_data_bits_7_14 = io_wgt_rd_data_bits_7_14; // @[TensorGemm.scala 346:19:@20857.4]
  assign mvc_io_wgt_data_bits_7_15 = io_wgt_rd_data_bits_7_15; // @[TensorGemm.scala 346:19:@20858.4]
  assign mvc_io_wgt_data_bits_8_0 = io_wgt_rd_data_bits_8_0; // @[TensorGemm.scala 346:19:@20859.4]
  assign mvc_io_wgt_data_bits_8_1 = io_wgt_rd_data_bits_8_1; // @[TensorGemm.scala 346:19:@20860.4]
  assign mvc_io_wgt_data_bits_8_2 = io_wgt_rd_data_bits_8_2; // @[TensorGemm.scala 346:19:@20861.4]
  assign mvc_io_wgt_data_bits_8_3 = io_wgt_rd_data_bits_8_3; // @[TensorGemm.scala 346:19:@20862.4]
  assign mvc_io_wgt_data_bits_8_4 = io_wgt_rd_data_bits_8_4; // @[TensorGemm.scala 346:19:@20863.4]
  assign mvc_io_wgt_data_bits_8_5 = io_wgt_rd_data_bits_8_5; // @[TensorGemm.scala 346:19:@20864.4]
  assign mvc_io_wgt_data_bits_8_6 = io_wgt_rd_data_bits_8_6; // @[TensorGemm.scala 346:19:@20865.4]
  assign mvc_io_wgt_data_bits_8_7 = io_wgt_rd_data_bits_8_7; // @[TensorGemm.scala 346:19:@20866.4]
  assign mvc_io_wgt_data_bits_8_8 = io_wgt_rd_data_bits_8_8; // @[TensorGemm.scala 346:19:@20867.4]
  assign mvc_io_wgt_data_bits_8_9 = io_wgt_rd_data_bits_8_9; // @[TensorGemm.scala 346:19:@20868.4]
  assign mvc_io_wgt_data_bits_8_10 = io_wgt_rd_data_bits_8_10; // @[TensorGemm.scala 346:19:@20869.4]
  assign mvc_io_wgt_data_bits_8_11 = io_wgt_rd_data_bits_8_11; // @[TensorGemm.scala 346:19:@20870.4]
  assign mvc_io_wgt_data_bits_8_12 = io_wgt_rd_data_bits_8_12; // @[TensorGemm.scala 346:19:@20871.4]
  assign mvc_io_wgt_data_bits_8_13 = io_wgt_rd_data_bits_8_13; // @[TensorGemm.scala 346:19:@20872.4]
  assign mvc_io_wgt_data_bits_8_14 = io_wgt_rd_data_bits_8_14; // @[TensorGemm.scala 346:19:@20873.4]
  assign mvc_io_wgt_data_bits_8_15 = io_wgt_rd_data_bits_8_15; // @[TensorGemm.scala 346:19:@20874.4]
  assign mvc_io_wgt_data_bits_9_0 = io_wgt_rd_data_bits_9_0; // @[TensorGemm.scala 346:19:@20875.4]
  assign mvc_io_wgt_data_bits_9_1 = io_wgt_rd_data_bits_9_1; // @[TensorGemm.scala 346:19:@20876.4]
  assign mvc_io_wgt_data_bits_9_2 = io_wgt_rd_data_bits_9_2; // @[TensorGemm.scala 346:19:@20877.4]
  assign mvc_io_wgt_data_bits_9_3 = io_wgt_rd_data_bits_9_3; // @[TensorGemm.scala 346:19:@20878.4]
  assign mvc_io_wgt_data_bits_9_4 = io_wgt_rd_data_bits_9_4; // @[TensorGemm.scala 346:19:@20879.4]
  assign mvc_io_wgt_data_bits_9_5 = io_wgt_rd_data_bits_9_5; // @[TensorGemm.scala 346:19:@20880.4]
  assign mvc_io_wgt_data_bits_9_6 = io_wgt_rd_data_bits_9_6; // @[TensorGemm.scala 346:19:@20881.4]
  assign mvc_io_wgt_data_bits_9_7 = io_wgt_rd_data_bits_9_7; // @[TensorGemm.scala 346:19:@20882.4]
  assign mvc_io_wgt_data_bits_9_8 = io_wgt_rd_data_bits_9_8; // @[TensorGemm.scala 346:19:@20883.4]
  assign mvc_io_wgt_data_bits_9_9 = io_wgt_rd_data_bits_9_9; // @[TensorGemm.scala 346:19:@20884.4]
  assign mvc_io_wgt_data_bits_9_10 = io_wgt_rd_data_bits_9_10; // @[TensorGemm.scala 346:19:@20885.4]
  assign mvc_io_wgt_data_bits_9_11 = io_wgt_rd_data_bits_9_11; // @[TensorGemm.scala 346:19:@20886.4]
  assign mvc_io_wgt_data_bits_9_12 = io_wgt_rd_data_bits_9_12; // @[TensorGemm.scala 346:19:@20887.4]
  assign mvc_io_wgt_data_bits_9_13 = io_wgt_rd_data_bits_9_13; // @[TensorGemm.scala 346:19:@20888.4]
  assign mvc_io_wgt_data_bits_9_14 = io_wgt_rd_data_bits_9_14; // @[TensorGemm.scala 346:19:@20889.4]
  assign mvc_io_wgt_data_bits_9_15 = io_wgt_rd_data_bits_9_15; // @[TensorGemm.scala 346:19:@20890.4]
  assign mvc_io_wgt_data_bits_10_0 = io_wgt_rd_data_bits_10_0; // @[TensorGemm.scala 346:19:@20891.4]
  assign mvc_io_wgt_data_bits_10_1 = io_wgt_rd_data_bits_10_1; // @[TensorGemm.scala 346:19:@20892.4]
  assign mvc_io_wgt_data_bits_10_2 = io_wgt_rd_data_bits_10_2; // @[TensorGemm.scala 346:19:@20893.4]
  assign mvc_io_wgt_data_bits_10_3 = io_wgt_rd_data_bits_10_3; // @[TensorGemm.scala 346:19:@20894.4]
  assign mvc_io_wgt_data_bits_10_4 = io_wgt_rd_data_bits_10_4; // @[TensorGemm.scala 346:19:@20895.4]
  assign mvc_io_wgt_data_bits_10_5 = io_wgt_rd_data_bits_10_5; // @[TensorGemm.scala 346:19:@20896.4]
  assign mvc_io_wgt_data_bits_10_6 = io_wgt_rd_data_bits_10_6; // @[TensorGemm.scala 346:19:@20897.4]
  assign mvc_io_wgt_data_bits_10_7 = io_wgt_rd_data_bits_10_7; // @[TensorGemm.scala 346:19:@20898.4]
  assign mvc_io_wgt_data_bits_10_8 = io_wgt_rd_data_bits_10_8; // @[TensorGemm.scala 346:19:@20899.4]
  assign mvc_io_wgt_data_bits_10_9 = io_wgt_rd_data_bits_10_9; // @[TensorGemm.scala 346:19:@20900.4]
  assign mvc_io_wgt_data_bits_10_10 = io_wgt_rd_data_bits_10_10; // @[TensorGemm.scala 346:19:@20901.4]
  assign mvc_io_wgt_data_bits_10_11 = io_wgt_rd_data_bits_10_11; // @[TensorGemm.scala 346:19:@20902.4]
  assign mvc_io_wgt_data_bits_10_12 = io_wgt_rd_data_bits_10_12; // @[TensorGemm.scala 346:19:@20903.4]
  assign mvc_io_wgt_data_bits_10_13 = io_wgt_rd_data_bits_10_13; // @[TensorGemm.scala 346:19:@20904.4]
  assign mvc_io_wgt_data_bits_10_14 = io_wgt_rd_data_bits_10_14; // @[TensorGemm.scala 346:19:@20905.4]
  assign mvc_io_wgt_data_bits_10_15 = io_wgt_rd_data_bits_10_15; // @[TensorGemm.scala 346:19:@20906.4]
  assign mvc_io_wgt_data_bits_11_0 = io_wgt_rd_data_bits_11_0; // @[TensorGemm.scala 346:19:@20907.4]
  assign mvc_io_wgt_data_bits_11_1 = io_wgt_rd_data_bits_11_1; // @[TensorGemm.scala 346:19:@20908.4]
  assign mvc_io_wgt_data_bits_11_2 = io_wgt_rd_data_bits_11_2; // @[TensorGemm.scala 346:19:@20909.4]
  assign mvc_io_wgt_data_bits_11_3 = io_wgt_rd_data_bits_11_3; // @[TensorGemm.scala 346:19:@20910.4]
  assign mvc_io_wgt_data_bits_11_4 = io_wgt_rd_data_bits_11_4; // @[TensorGemm.scala 346:19:@20911.4]
  assign mvc_io_wgt_data_bits_11_5 = io_wgt_rd_data_bits_11_5; // @[TensorGemm.scala 346:19:@20912.4]
  assign mvc_io_wgt_data_bits_11_6 = io_wgt_rd_data_bits_11_6; // @[TensorGemm.scala 346:19:@20913.4]
  assign mvc_io_wgt_data_bits_11_7 = io_wgt_rd_data_bits_11_7; // @[TensorGemm.scala 346:19:@20914.4]
  assign mvc_io_wgt_data_bits_11_8 = io_wgt_rd_data_bits_11_8; // @[TensorGemm.scala 346:19:@20915.4]
  assign mvc_io_wgt_data_bits_11_9 = io_wgt_rd_data_bits_11_9; // @[TensorGemm.scala 346:19:@20916.4]
  assign mvc_io_wgt_data_bits_11_10 = io_wgt_rd_data_bits_11_10; // @[TensorGemm.scala 346:19:@20917.4]
  assign mvc_io_wgt_data_bits_11_11 = io_wgt_rd_data_bits_11_11; // @[TensorGemm.scala 346:19:@20918.4]
  assign mvc_io_wgt_data_bits_11_12 = io_wgt_rd_data_bits_11_12; // @[TensorGemm.scala 346:19:@20919.4]
  assign mvc_io_wgt_data_bits_11_13 = io_wgt_rd_data_bits_11_13; // @[TensorGemm.scala 346:19:@20920.4]
  assign mvc_io_wgt_data_bits_11_14 = io_wgt_rd_data_bits_11_14; // @[TensorGemm.scala 346:19:@20921.4]
  assign mvc_io_wgt_data_bits_11_15 = io_wgt_rd_data_bits_11_15; // @[TensorGemm.scala 346:19:@20922.4]
  assign mvc_io_wgt_data_bits_12_0 = io_wgt_rd_data_bits_12_0; // @[TensorGemm.scala 346:19:@20923.4]
  assign mvc_io_wgt_data_bits_12_1 = io_wgt_rd_data_bits_12_1; // @[TensorGemm.scala 346:19:@20924.4]
  assign mvc_io_wgt_data_bits_12_2 = io_wgt_rd_data_bits_12_2; // @[TensorGemm.scala 346:19:@20925.4]
  assign mvc_io_wgt_data_bits_12_3 = io_wgt_rd_data_bits_12_3; // @[TensorGemm.scala 346:19:@20926.4]
  assign mvc_io_wgt_data_bits_12_4 = io_wgt_rd_data_bits_12_4; // @[TensorGemm.scala 346:19:@20927.4]
  assign mvc_io_wgt_data_bits_12_5 = io_wgt_rd_data_bits_12_5; // @[TensorGemm.scala 346:19:@20928.4]
  assign mvc_io_wgt_data_bits_12_6 = io_wgt_rd_data_bits_12_6; // @[TensorGemm.scala 346:19:@20929.4]
  assign mvc_io_wgt_data_bits_12_7 = io_wgt_rd_data_bits_12_7; // @[TensorGemm.scala 346:19:@20930.4]
  assign mvc_io_wgt_data_bits_12_8 = io_wgt_rd_data_bits_12_8; // @[TensorGemm.scala 346:19:@20931.4]
  assign mvc_io_wgt_data_bits_12_9 = io_wgt_rd_data_bits_12_9; // @[TensorGemm.scala 346:19:@20932.4]
  assign mvc_io_wgt_data_bits_12_10 = io_wgt_rd_data_bits_12_10; // @[TensorGemm.scala 346:19:@20933.4]
  assign mvc_io_wgt_data_bits_12_11 = io_wgt_rd_data_bits_12_11; // @[TensorGemm.scala 346:19:@20934.4]
  assign mvc_io_wgt_data_bits_12_12 = io_wgt_rd_data_bits_12_12; // @[TensorGemm.scala 346:19:@20935.4]
  assign mvc_io_wgt_data_bits_12_13 = io_wgt_rd_data_bits_12_13; // @[TensorGemm.scala 346:19:@20936.4]
  assign mvc_io_wgt_data_bits_12_14 = io_wgt_rd_data_bits_12_14; // @[TensorGemm.scala 346:19:@20937.4]
  assign mvc_io_wgt_data_bits_12_15 = io_wgt_rd_data_bits_12_15; // @[TensorGemm.scala 346:19:@20938.4]
  assign mvc_io_wgt_data_bits_13_0 = io_wgt_rd_data_bits_13_0; // @[TensorGemm.scala 346:19:@20939.4]
  assign mvc_io_wgt_data_bits_13_1 = io_wgt_rd_data_bits_13_1; // @[TensorGemm.scala 346:19:@20940.4]
  assign mvc_io_wgt_data_bits_13_2 = io_wgt_rd_data_bits_13_2; // @[TensorGemm.scala 346:19:@20941.4]
  assign mvc_io_wgt_data_bits_13_3 = io_wgt_rd_data_bits_13_3; // @[TensorGemm.scala 346:19:@20942.4]
  assign mvc_io_wgt_data_bits_13_4 = io_wgt_rd_data_bits_13_4; // @[TensorGemm.scala 346:19:@20943.4]
  assign mvc_io_wgt_data_bits_13_5 = io_wgt_rd_data_bits_13_5; // @[TensorGemm.scala 346:19:@20944.4]
  assign mvc_io_wgt_data_bits_13_6 = io_wgt_rd_data_bits_13_6; // @[TensorGemm.scala 346:19:@20945.4]
  assign mvc_io_wgt_data_bits_13_7 = io_wgt_rd_data_bits_13_7; // @[TensorGemm.scala 346:19:@20946.4]
  assign mvc_io_wgt_data_bits_13_8 = io_wgt_rd_data_bits_13_8; // @[TensorGemm.scala 346:19:@20947.4]
  assign mvc_io_wgt_data_bits_13_9 = io_wgt_rd_data_bits_13_9; // @[TensorGemm.scala 346:19:@20948.4]
  assign mvc_io_wgt_data_bits_13_10 = io_wgt_rd_data_bits_13_10; // @[TensorGemm.scala 346:19:@20949.4]
  assign mvc_io_wgt_data_bits_13_11 = io_wgt_rd_data_bits_13_11; // @[TensorGemm.scala 346:19:@20950.4]
  assign mvc_io_wgt_data_bits_13_12 = io_wgt_rd_data_bits_13_12; // @[TensorGemm.scala 346:19:@20951.4]
  assign mvc_io_wgt_data_bits_13_13 = io_wgt_rd_data_bits_13_13; // @[TensorGemm.scala 346:19:@20952.4]
  assign mvc_io_wgt_data_bits_13_14 = io_wgt_rd_data_bits_13_14; // @[TensorGemm.scala 346:19:@20953.4]
  assign mvc_io_wgt_data_bits_13_15 = io_wgt_rd_data_bits_13_15; // @[TensorGemm.scala 346:19:@20954.4]
  assign mvc_io_wgt_data_bits_14_0 = io_wgt_rd_data_bits_14_0; // @[TensorGemm.scala 346:19:@20955.4]
  assign mvc_io_wgt_data_bits_14_1 = io_wgt_rd_data_bits_14_1; // @[TensorGemm.scala 346:19:@20956.4]
  assign mvc_io_wgt_data_bits_14_2 = io_wgt_rd_data_bits_14_2; // @[TensorGemm.scala 346:19:@20957.4]
  assign mvc_io_wgt_data_bits_14_3 = io_wgt_rd_data_bits_14_3; // @[TensorGemm.scala 346:19:@20958.4]
  assign mvc_io_wgt_data_bits_14_4 = io_wgt_rd_data_bits_14_4; // @[TensorGemm.scala 346:19:@20959.4]
  assign mvc_io_wgt_data_bits_14_5 = io_wgt_rd_data_bits_14_5; // @[TensorGemm.scala 346:19:@20960.4]
  assign mvc_io_wgt_data_bits_14_6 = io_wgt_rd_data_bits_14_6; // @[TensorGemm.scala 346:19:@20961.4]
  assign mvc_io_wgt_data_bits_14_7 = io_wgt_rd_data_bits_14_7; // @[TensorGemm.scala 346:19:@20962.4]
  assign mvc_io_wgt_data_bits_14_8 = io_wgt_rd_data_bits_14_8; // @[TensorGemm.scala 346:19:@20963.4]
  assign mvc_io_wgt_data_bits_14_9 = io_wgt_rd_data_bits_14_9; // @[TensorGemm.scala 346:19:@20964.4]
  assign mvc_io_wgt_data_bits_14_10 = io_wgt_rd_data_bits_14_10; // @[TensorGemm.scala 346:19:@20965.4]
  assign mvc_io_wgt_data_bits_14_11 = io_wgt_rd_data_bits_14_11; // @[TensorGemm.scala 346:19:@20966.4]
  assign mvc_io_wgt_data_bits_14_12 = io_wgt_rd_data_bits_14_12; // @[TensorGemm.scala 346:19:@20967.4]
  assign mvc_io_wgt_data_bits_14_13 = io_wgt_rd_data_bits_14_13; // @[TensorGemm.scala 346:19:@20968.4]
  assign mvc_io_wgt_data_bits_14_14 = io_wgt_rd_data_bits_14_14; // @[TensorGemm.scala 346:19:@20969.4]
  assign mvc_io_wgt_data_bits_14_15 = io_wgt_rd_data_bits_14_15; // @[TensorGemm.scala 346:19:@20970.4]
  assign mvc_io_wgt_data_bits_15_0 = io_wgt_rd_data_bits_15_0; // @[TensorGemm.scala 346:19:@20971.4]
  assign mvc_io_wgt_data_bits_15_1 = io_wgt_rd_data_bits_15_1; // @[TensorGemm.scala 346:19:@20972.4]
  assign mvc_io_wgt_data_bits_15_2 = io_wgt_rd_data_bits_15_2; // @[TensorGemm.scala 346:19:@20973.4]
  assign mvc_io_wgt_data_bits_15_3 = io_wgt_rd_data_bits_15_3; // @[TensorGemm.scala 346:19:@20974.4]
  assign mvc_io_wgt_data_bits_15_4 = io_wgt_rd_data_bits_15_4; // @[TensorGemm.scala 346:19:@20975.4]
  assign mvc_io_wgt_data_bits_15_5 = io_wgt_rd_data_bits_15_5; // @[TensorGemm.scala 346:19:@20976.4]
  assign mvc_io_wgt_data_bits_15_6 = io_wgt_rd_data_bits_15_6; // @[TensorGemm.scala 346:19:@20977.4]
  assign mvc_io_wgt_data_bits_15_7 = io_wgt_rd_data_bits_15_7; // @[TensorGemm.scala 346:19:@20978.4]
  assign mvc_io_wgt_data_bits_15_8 = io_wgt_rd_data_bits_15_8; // @[TensorGemm.scala 346:19:@20979.4]
  assign mvc_io_wgt_data_bits_15_9 = io_wgt_rd_data_bits_15_9; // @[TensorGemm.scala 346:19:@20980.4]
  assign mvc_io_wgt_data_bits_15_10 = io_wgt_rd_data_bits_15_10; // @[TensorGemm.scala 346:19:@20981.4]
  assign mvc_io_wgt_data_bits_15_11 = io_wgt_rd_data_bits_15_11; // @[TensorGemm.scala 346:19:@20982.4]
  assign mvc_io_wgt_data_bits_15_12 = io_wgt_rd_data_bits_15_12; // @[TensorGemm.scala 346:19:@20983.4]
  assign mvc_io_wgt_data_bits_15_13 = io_wgt_rd_data_bits_15_13; // @[TensorGemm.scala 346:19:@20984.4]
  assign mvc_io_wgt_data_bits_15_14 = io_wgt_rd_data_bits_15_14; // @[TensorGemm.scala 346:19:@20985.4]
  assign mvc_io_wgt_data_bits_15_15 = io_wgt_rd_data_bits_15_15; // @[TensorGemm.scala 346:19:@20986.4]
  assign mvc_io_acc_i_data_valid = io_acc_rd_data_valid; // @[TensorGemm.scala 347:21:@21004.4]
  assign mvc_io_acc_i_data_bits_0_0 = io_acc_rd_data_bits_0_0; // @[TensorGemm.scala 347:21:@20988.4]
  assign mvc_io_acc_i_data_bits_0_1 = io_acc_rd_data_bits_0_1; // @[TensorGemm.scala 347:21:@20989.4]
  assign mvc_io_acc_i_data_bits_0_2 = io_acc_rd_data_bits_0_2; // @[TensorGemm.scala 347:21:@20990.4]
  assign mvc_io_acc_i_data_bits_0_3 = io_acc_rd_data_bits_0_3; // @[TensorGemm.scala 347:21:@20991.4]
  assign mvc_io_acc_i_data_bits_0_4 = io_acc_rd_data_bits_0_4; // @[TensorGemm.scala 347:21:@20992.4]
  assign mvc_io_acc_i_data_bits_0_5 = io_acc_rd_data_bits_0_5; // @[TensorGemm.scala 347:21:@20993.4]
  assign mvc_io_acc_i_data_bits_0_6 = io_acc_rd_data_bits_0_6; // @[TensorGemm.scala 347:21:@20994.4]
  assign mvc_io_acc_i_data_bits_0_7 = io_acc_rd_data_bits_0_7; // @[TensorGemm.scala 347:21:@20995.4]
  assign mvc_io_acc_i_data_bits_0_8 = io_acc_rd_data_bits_0_8; // @[TensorGemm.scala 347:21:@20996.4]
  assign mvc_io_acc_i_data_bits_0_9 = io_acc_rd_data_bits_0_9; // @[TensorGemm.scala 347:21:@20997.4]
  assign mvc_io_acc_i_data_bits_0_10 = io_acc_rd_data_bits_0_10; // @[TensorGemm.scala 347:21:@20998.4]
  assign mvc_io_acc_i_data_bits_0_11 = io_acc_rd_data_bits_0_11; // @[TensorGemm.scala 347:21:@20999.4]
  assign mvc_io_acc_i_data_bits_0_12 = io_acc_rd_data_bits_0_12; // @[TensorGemm.scala 347:21:@21000.4]
  assign mvc_io_acc_i_data_bits_0_13 = io_acc_rd_data_bits_0_13; // @[TensorGemm.scala 347:21:@21001.4]
  assign mvc_io_acc_i_data_bits_0_14 = io_acc_rd_data_bits_0_14; // @[TensorGemm.scala 347:21:@21002.4]
  assign mvc_io_acc_i_data_bits_0_15 = io_acc_rd_data_bits_0_15; // @[TensorGemm.scala 347:21:@21003.4]
  assign wrpipe_clock = clock; // @[:@20204.4]
  assign wrpipe_reset = reset; // @[:@20205.4]
  assign wrpipe_io_enq_valid = _T_7689 & _T_7830; // @[TensorGemm.scala 322:23:@20421.4]
  assign wrpipe_io_enq_bits = uop_acc; // @[TensorGemm.scala 323:22:@20422.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  uop_idx = _RAND_1[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  uop_acc = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  uop_inp = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  uop_wgt = _RAND_4[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  cnt_o = _RAND_5[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  acc_o = _RAND_6[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inp_o = _RAND_7[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wgt_o = _RAND_8[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  cnt_i = _RAND_9[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  acc_i = _RAND_10[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  inp_i = _RAND_11[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wgt_i = _RAND_12[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_7713) begin
        if (io_start) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_7714) begin
          state <= 3'h2;
        end else begin
          if (_T_7715) begin
            state <= 3'h3;
          end else begin
            if (_T_7716) begin
              state <= 3'h4;
            end else begin
              if (_T_7717) begin
                if (_T_7734) begin
                  if (_T_7736) begin
                    state <= 3'h5;
                  end else begin
                    state <= 3'h0;
                  end
                end else begin
                  state <= 3'h1;
                end
              end else begin
                if (_T_7737) begin
                  if (_T_7688) begin
                    state <= 3'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_7762) begin
      uop_idx <= {{1'd0}, dec_uop_begin};
    end else begin
      if (_T_7765) begin
        uop_idx <= _T_7768;
      end
    end
    if (_T_7822) begin
      uop_acc <= _T_7824;
    end
    if (_T_7822) begin
      uop_inp <= _T_7826;
    end
    if (_T_7822) begin
      uop_wgt <= _T_7828;
    end
    if (_T_7740) begin
      cnt_o <= 14'h0;
    end else begin
      if (_T_7786) begin
        cnt_o <= _T_7789;
      end
    end
    if (_T_7740) begin
      acc_o <= 14'h0;
    end else begin
      if (_T_7786) begin
        acc_o <= _T_7791;
      end
    end
    if (_T_7740) begin
      inp_o <= 14'h0;
    end else begin
      if (_T_7786) begin
        inp_o <= _T_7793;
      end
    end
    if (_T_7740) begin
      wgt_o <= 14'h0;
    end else begin
      if (_T_7786) begin
        wgt_o <= _T_7795;
      end
    end
    if (_T_7740) begin
      cnt_i <= 14'h0;
    end else begin
      if (_T_7803) begin
        cnt_i <= 14'h0;
      end else begin
        if (_T_7761) begin
          cnt_i <= _T_7814;
        end
      end
    end
    if (_T_7740) begin
      acc_i <= 14'h0;
    end else begin
      if (_T_7803) begin
        acc_i <= acc_o;
      end else begin
        if (_T_7761) begin
          acc_i <= _T_7816;
        end
      end
    end
    if (_T_7740) begin
      inp_i <= 14'h0;
    end else begin
      if (_T_7803) begin
        inp_i <= inp_o;
      end else begin
        if (_T_7761) begin
          inp_i <= _T_7818;
        end
      end
    end
    if (_T_7740) begin
      wgt_i <= 14'h0;
    end else begin
      if (_T_7803) begin
        wgt_i <= wgt_o;
      end else begin
        if (_T_7761) begin
          wgt_i <= _T_7820;
        end
      end
    end
    if (_T_7740) begin
      inflight <= 5'h0;
    end else begin
      if (_T_7743) begin
        if (!(_T_7745)) begin
          if (_T_7744) begin
            inflight <= _T_7749;
          end else begin
            if (mvc_io_acc_o_data_valid) begin
              inflight <= _T_7753;
            end
          end
        end
      end
    end
  end
endmodule
module Alu( // @[:@21049.2]
  input  [2:0]  io_opcode, // @[:@21052.4]
  input  [31:0] io_a, // @[:@21052.4]
  input  [31:0] io_b, // @[:@21052.4]
  output [31:0] io_y // @[:@21052.4]
);
  wire [31:0] ub; // @[TensorAlu.scala 37:17:@21054.4]
  wire [4:0] _T_13; // @[TensorAlu.scala 39:14:@21055.4]
  wire [4:0] _T_14; // @[TensorAlu.scala 39:11:@21056.4]
  wire [5:0] _T_16; // @[TensorAlu.scala 39:29:@21057.4]
  wire [4:0] m; // @[TensorAlu.scala 39:29:@21058.4]
  wire  _T_17; // @[TensorAlu.scala 42:26:@21060.4]
  wire [31:0] fop_0; // @[TensorAlu.scala 42:20:@21061.4]
  wire [31:0] fop_1; // @[TensorAlu.scala 42:50:@21063.4]
  wire [32:0] _T_19; // @[TensorAlu.scala 43:10:@21064.4]
  wire [31:0] _T_20; // @[TensorAlu.scala 43:10:@21065.4]
  wire [31:0] fop_2; // @[TensorAlu.scala 43:10:@21066.4]
  wire [31:0] fop_3; // @[TensorAlu.scala 43:23:@21067.4]
  wire [62:0] _GEN_0; // @[TensorAlu.scala 43:34:@21068.4]
  wire [62:0] fop_4; // @[TensorAlu.scala 43:34:@21068.4]
  wire  _T_21; // @[Mux.scala 46:19:@21069.4]
  wire [62:0] _T_22; // @[Mux.scala 46:16:@21070.4]
  wire  _T_23; // @[Mux.scala 46:19:@21071.4]
  wire [62:0] _T_24; // @[Mux.scala 46:16:@21072.4]
  wire  _T_25; // @[Mux.scala 46:19:@21073.4]
  wire [62:0] _T_26; // @[Mux.scala 46:16:@21074.4]
  wire  _T_27; // @[Mux.scala 46:19:@21075.4]
  wire [62:0] _T_28; // @[Mux.scala 46:16:@21076.4]
  wire  _T_29; // @[Mux.scala 46:19:@21077.4]
  wire [62:0] _T_30; // @[Mux.scala 46:16:@21078.4]
  wire [31:0] _GEN_1; // @[TensorAlu.scala 46:8:@21079.4]
  assign ub = $unsigned(io_b); // @[TensorAlu.scala 37:17:@21054.4]
  assign _T_13 = ub[4:0]; // @[TensorAlu.scala 39:14:@21055.4]
  assign _T_14 = ~ _T_13; // @[TensorAlu.scala 39:11:@21056.4]
  assign _T_16 = _T_14 + 5'h1; // @[TensorAlu.scala 39:29:@21057.4]
  assign m = _T_14 + 5'h1; // @[TensorAlu.scala 39:29:@21058.4]
  assign _T_17 = $signed(io_a) < $signed(io_b); // @[TensorAlu.scala 42:26:@21060.4]
  assign fop_0 = _T_17 ? $signed(io_a) : $signed(io_b); // @[TensorAlu.scala 42:20:@21061.4]
  assign fop_1 = _T_17 ? $signed(io_b) : $signed(io_a); // @[TensorAlu.scala 42:50:@21063.4]
  assign _T_19 = $signed(io_a) + $signed(io_b); // @[TensorAlu.scala 43:10:@21064.4]
  assign _T_20 = $signed(io_a) + $signed(io_b); // @[TensorAlu.scala 43:10:@21065.4]
  assign fop_2 = $signed(_T_20); // @[TensorAlu.scala 43:10:@21066.4]
  assign fop_3 = $signed(io_a) >>> _T_13; // @[TensorAlu.scala 43:23:@21067.4]
  assign _GEN_0 = {{31{io_a[31]}},io_a}; // @[TensorAlu.scala 43:34:@21068.4]
  assign fop_4 = $signed(_GEN_0) << m; // @[TensorAlu.scala 43:34:@21068.4]
  assign _T_21 = 3'h4 == io_opcode; // @[Mux.scala 46:19:@21069.4]
  assign _T_22 = _T_21 ? $signed(fop_4) : $signed({{31{io_a[31]}},io_a}); // @[Mux.scala 46:16:@21070.4]
  assign _T_23 = 3'h3 == io_opcode; // @[Mux.scala 46:19:@21071.4]
  assign _T_24 = _T_23 ? $signed({{31{fop_3[31]}},fop_3}) : $signed(_T_22); // @[Mux.scala 46:16:@21072.4]
  assign _T_25 = 3'h2 == io_opcode; // @[Mux.scala 46:19:@21073.4]
  assign _T_26 = _T_25 ? $signed({{31{fop_2[31]}},fop_2}) : $signed(_T_24); // @[Mux.scala 46:16:@21074.4]
  assign _T_27 = 3'h1 == io_opcode; // @[Mux.scala 46:19:@21075.4]
  assign _T_28 = _T_27 ? $signed({{31{fop_1[31]}},fop_1}) : $signed(_T_26); // @[Mux.scala 46:16:@21076.4]
  assign _T_29 = 3'h0 == io_opcode; // @[Mux.scala 46:19:@21077.4]
  assign _T_30 = _T_29 ? $signed({{31{fop_0[31]}},fop_0}) : $signed(_T_28); // @[Mux.scala 46:16:@21078.4]
  assign _GEN_1 = _T_30[31:0]; // @[TensorAlu.scala 46:8:@21079.4]
  assign io_y = $signed(_GEN_1); // @[TensorAlu.scala 46:8:@21079.4]
endmodule
module AluReg( // @[:@21081.2]
  input         clock, // @[:@21082.4]
  input  [2:0]  io_opcode, // @[:@21084.4]
  input         io_a_valid, // @[:@21084.4]
  input  [31:0] io_a_bits, // @[:@21084.4]
  input         io_b_valid, // @[:@21084.4]
  input  [31:0] io_b_bits, // @[:@21084.4]
  output        io_y_valid, // @[:@21084.4]
  output [31:0] io_y_bits // @[:@21084.4]
);
  wire [2:0] alu_io_opcode; // @[TensorAlu.scala 57:19:@21086.4]
  wire [31:0] alu_io_a; // @[TensorAlu.scala 57:19:@21086.4]
  wire [31:0] alu_io_b; // @[TensorAlu.scala 57:19:@21086.4]
  wire [31:0] alu_io_y; // @[TensorAlu.scala 57:19:@21086.4]
  reg [31:0] rA; // @[Reg.scala 11:16:@21089.4]
  reg [31:0] _RAND_0;
  reg [31:0] rB; // @[Reg.scala 11:16:@21093.4]
  reg [31:0] _RAND_1;
  reg  valid; // @[TensorAlu.scala 60:22:@21097.4]
  reg [31:0] _RAND_2;
  Alu alu ( // @[TensorAlu.scala 57:19:@21086.4]
    .io_opcode(alu_io_opcode),
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_y(alu_io_y)
  );
  assign io_y_valid = valid; // @[TensorAlu.scala 69:14:@21104.4]
  assign io_y_bits = $unsigned(alu_io_y); // @[TensorAlu.scala 70:13:@21106.4]
  assign alu_io_opcode = io_opcode; // @[TensorAlu.scala 62:17:@21099.4]
  assign alu_io_a = $signed(rA); // @[TensorAlu.scala 65:12:@21101.4]
  assign alu_io_b = $signed(rB); // @[TensorAlu.scala 66:12:@21103.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rA = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rB = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_a_valid) begin
      rA <= io_a_bits;
    end
    if (io_b_valid) begin
      rB <= io_b_bits;
    end
    valid <= io_b_valid;
  end
endmodule
module AluVector( // @[:@21993.2]
  input         clock, // @[:@21994.4]
  input  [2:0]  io_opcode, // @[:@21996.4]
  input         io_acc_a_data_valid, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_0, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_1, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_2, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_3, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_4, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_5, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_6, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_7, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_8, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_9, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_10, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_11, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_12, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_13, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_14, // @[:@21996.4]
  input  [31:0] io_acc_a_data_bits_0_15, // @[:@21996.4]
  input         io_acc_b_data_valid, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_0, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_1, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_2, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_3, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_4, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_5, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_6, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_7, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_8, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_9, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_10, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_11, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_12, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_13, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_14, // @[:@21996.4]
  input  [31:0] io_acc_b_data_bits_0_15, // @[:@21996.4]
  output        io_acc_y_data_valid, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_0, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_1, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_2, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_3, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_4, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_5, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_6, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_7, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_8, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_9, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_10, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_11, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_12, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_13, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_14, // @[:@21996.4]
  output [31:0] io_acc_y_data_bits_0_15, // @[:@21996.4]
  output        io_out_data_valid, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_0, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_1, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_2, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_3, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_4, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_5, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_6, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_7, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_8, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_9, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_10, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_11, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_12, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_13, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_14, // @[:@21996.4]
  output [7:0]  io_out_data_bits_0_15 // @[:@21996.4]
);
  wire  f_0_clock; // @[TensorAlu.scala 83:36:@21998.4]
  wire [2:0] f_0_io_opcode; // @[TensorAlu.scala 83:36:@21998.4]
  wire  f_0_io_a_valid; // @[TensorAlu.scala 83:36:@21998.4]
  wire [31:0] f_0_io_a_bits; // @[TensorAlu.scala 83:36:@21998.4]
  wire  f_0_io_b_valid; // @[TensorAlu.scala 83:36:@21998.4]
  wire [31:0] f_0_io_b_bits; // @[TensorAlu.scala 83:36:@21998.4]
  wire  f_0_io_y_valid; // @[TensorAlu.scala 83:36:@21998.4]
  wire [31:0] f_0_io_y_bits; // @[TensorAlu.scala 83:36:@21998.4]
  wire  f_1_clock; // @[TensorAlu.scala 83:36:@22001.4]
  wire [2:0] f_1_io_opcode; // @[TensorAlu.scala 83:36:@22001.4]
  wire  f_1_io_a_valid; // @[TensorAlu.scala 83:36:@22001.4]
  wire [31:0] f_1_io_a_bits; // @[TensorAlu.scala 83:36:@22001.4]
  wire  f_1_io_b_valid; // @[TensorAlu.scala 83:36:@22001.4]
  wire [31:0] f_1_io_b_bits; // @[TensorAlu.scala 83:36:@22001.4]
  wire  f_1_io_y_valid; // @[TensorAlu.scala 83:36:@22001.4]
  wire [31:0] f_1_io_y_bits; // @[TensorAlu.scala 83:36:@22001.4]
  wire  f_2_clock; // @[TensorAlu.scala 83:36:@22004.4]
  wire [2:0] f_2_io_opcode; // @[TensorAlu.scala 83:36:@22004.4]
  wire  f_2_io_a_valid; // @[TensorAlu.scala 83:36:@22004.4]
  wire [31:0] f_2_io_a_bits; // @[TensorAlu.scala 83:36:@22004.4]
  wire  f_2_io_b_valid; // @[TensorAlu.scala 83:36:@22004.4]
  wire [31:0] f_2_io_b_bits; // @[TensorAlu.scala 83:36:@22004.4]
  wire  f_2_io_y_valid; // @[TensorAlu.scala 83:36:@22004.4]
  wire [31:0] f_2_io_y_bits; // @[TensorAlu.scala 83:36:@22004.4]
  wire  f_3_clock; // @[TensorAlu.scala 83:36:@22007.4]
  wire [2:0] f_3_io_opcode; // @[TensorAlu.scala 83:36:@22007.4]
  wire  f_3_io_a_valid; // @[TensorAlu.scala 83:36:@22007.4]
  wire [31:0] f_3_io_a_bits; // @[TensorAlu.scala 83:36:@22007.4]
  wire  f_3_io_b_valid; // @[TensorAlu.scala 83:36:@22007.4]
  wire [31:0] f_3_io_b_bits; // @[TensorAlu.scala 83:36:@22007.4]
  wire  f_3_io_y_valid; // @[TensorAlu.scala 83:36:@22007.4]
  wire [31:0] f_3_io_y_bits; // @[TensorAlu.scala 83:36:@22007.4]
  wire  f_4_clock; // @[TensorAlu.scala 83:36:@22010.4]
  wire [2:0] f_4_io_opcode; // @[TensorAlu.scala 83:36:@22010.4]
  wire  f_4_io_a_valid; // @[TensorAlu.scala 83:36:@22010.4]
  wire [31:0] f_4_io_a_bits; // @[TensorAlu.scala 83:36:@22010.4]
  wire  f_4_io_b_valid; // @[TensorAlu.scala 83:36:@22010.4]
  wire [31:0] f_4_io_b_bits; // @[TensorAlu.scala 83:36:@22010.4]
  wire  f_4_io_y_valid; // @[TensorAlu.scala 83:36:@22010.4]
  wire [31:0] f_4_io_y_bits; // @[TensorAlu.scala 83:36:@22010.4]
  wire  f_5_clock; // @[TensorAlu.scala 83:36:@22013.4]
  wire [2:0] f_5_io_opcode; // @[TensorAlu.scala 83:36:@22013.4]
  wire  f_5_io_a_valid; // @[TensorAlu.scala 83:36:@22013.4]
  wire [31:0] f_5_io_a_bits; // @[TensorAlu.scala 83:36:@22013.4]
  wire  f_5_io_b_valid; // @[TensorAlu.scala 83:36:@22013.4]
  wire [31:0] f_5_io_b_bits; // @[TensorAlu.scala 83:36:@22013.4]
  wire  f_5_io_y_valid; // @[TensorAlu.scala 83:36:@22013.4]
  wire [31:0] f_5_io_y_bits; // @[TensorAlu.scala 83:36:@22013.4]
  wire  f_6_clock; // @[TensorAlu.scala 83:36:@22016.4]
  wire [2:0] f_6_io_opcode; // @[TensorAlu.scala 83:36:@22016.4]
  wire  f_6_io_a_valid; // @[TensorAlu.scala 83:36:@22016.4]
  wire [31:0] f_6_io_a_bits; // @[TensorAlu.scala 83:36:@22016.4]
  wire  f_6_io_b_valid; // @[TensorAlu.scala 83:36:@22016.4]
  wire [31:0] f_6_io_b_bits; // @[TensorAlu.scala 83:36:@22016.4]
  wire  f_6_io_y_valid; // @[TensorAlu.scala 83:36:@22016.4]
  wire [31:0] f_6_io_y_bits; // @[TensorAlu.scala 83:36:@22016.4]
  wire  f_7_clock; // @[TensorAlu.scala 83:36:@22019.4]
  wire [2:0] f_7_io_opcode; // @[TensorAlu.scala 83:36:@22019.4]
  wire  f_7_io_a_valid; // @[TensorAlu.scala 83:36:@22019.4]
  wire [31:0] f_7_io_a_bits; // @[TensorAlu.scala 83:36:@22019.4]
  wire  f_7_io_b_valid; // @[TensorAlu.scala 83:36:@22019.4]
  wire [31:0] f_7_io_b_bits; // @[TensorAlu.scala 83:36:@22019.4]
  wire  f_7_io_y_valid; // @[TensorAlu.scala 83:36:@22019.4]
  wire [31:0] f_7_io_y_bits; // @[TensorAlu.scala 83:36:@22019.4]
  wire  f_8_clock; // @[TensorAlu.scala 83:36:@22022.4]
  wire [2:0] f_8_io_opcode; // @[TensorAlu.scala 83:36:@22022.4]
  wire  f_8_io_a_valid; // @[TensorAlu.scala 83:36:@22022.4]
  wire [31:0] f_8_io_a_bits; // @[TensorAlu.scala 83:36:@22022.4]
  wire  f_8_io_b_valid; // @[TensorAlu.scala 83:36:@22022.4]
  wire [31:0] f_8_io_b_bits; // @[TensorAlu.scala 83:36:@22022.4]
  wire  f_8_io_y_valid; // @[TensorAlu.scala 83:36:@22022.4]
  wire [31:0] f_8_io_y_bits; // @[TensorAlu.scala 83:36:@22022.4]
  wire  f_9_clock; // @[TensorAlu.scala 83:36:@22025.4]
  wire [2:0] f_9_io_opcode; // @[TensorAlu.scala 83:36:@22025.4]
  wire  f_9_io_a_valid; // @[TensorAlu.scala 83:36:@22025.4]
  wire [31:0] f_9_io_a_bits; // @[TensorAlu.scala 83:36:@22025.4]
  wire  f_9_io_b_valid; // @[TensorAlu.scala 83:36:@22025.4]
  wire [31:0] f_9_io_b_bits; // @[TensorAlu.scala 83:36:@22025.4]
  wire  f_9_io_y_valid; // @[TensorAlu.scala 83:36:@22025.4]
  wire [31:0] f_9_io_y_bits; // @[TensorAlu.scala 83:36:@22025.4]
  wire  f_10_clock; // @[TensorAlu.scala 83:36:@22028.4]
  wire [2:0] f_10_io_opcode; // @[TensorAlu.scala 83:36:@22028.4]
  wire  f_10_io_a_valid; // @[TensorAlu.scala 83:36:@22028.4]
  wire [31:0] f_10_io_a_bits; // @[TensorAlu.scala 83:36:@22028.4]
  wire  f_10_io_b_valid; // @[TensorAlu.scala 83:36:@22028.4]
  wire [31:0] f_10_io_b_bits; // @[TensorAlu.scala 83:36:@22028.4]
  wire  f_10_io_y_valid; // @[TensorAlu.scala 83:36:@22028.4]
  wire [31:0] f_10_io_y_bits; // @[TensorAlu.scala 83:36:@22028.4]
  wire  f_11_clock; // @[TensorAlu.scala 83:36:@22031.4]
  wire [2:0] f_11_io_opcode; // @[TensorAlu.scala 83:36:@22031.4]
  wire  f_11_io_a_valid; // @[TensorAlu.scala 83:36:@22031.4]
  wire [31:0] f_11_io_a_bits; // @[TensorAlu.scala 83:36:@22031.4]
  wire  f_11_io_b_valid; // @[TensorAlu.scala 83:36:@22031.4]
  wire [31:0] f_11_io_b_bits; // @[TensorAlu.scala 83:36:@22031.4]
  wire  f_11_io_y_valid; // @[TensorAlu.scala 83:36:@22031.4]
  wire [31:0] f_11_io_y_bits; // @[TensorAlu.scala 83:36:@22031.4]
  wire  f_12_clock; // @[TensorAlu.scala 83:36:@22034.4]
  wire [2:0] f_12_io_opcode; // @[TensorAlu.scala 83:36:@22034.4]
  wire  f_12_io_a_valid; // @[TensorAlu.scala 83:36:@22034.4]
  wire [31:0] f_12_io_a_bits; // @[TensorAlu.scala 83:36:@22034.4]
  wire  f_12_io_b_valid; // @[TensorAlu.scala 83:36:@22034.4]
  wire [31:0] f_12_io_b_bits; // @[TensorAlu.scala 83:36:@22034.4]
  wire  f_12_io_y_valid; // @[TensorAlu.scala 83:36:@22034.4]
  wire [31:0] f_12_io_y_bits; // @[TensorAlu.scala 83:36:@22034.4]
  wire  f_13_clock; // @[TensorAlu.scala 83:36:@22037.4]
  wire [2:0] f_13_io_opcode; // @[TensorAlu.scala 83:36:@22037.4]
  wire  f_13_io_a_valid; // @[TensorAlu.scala 83:36:@22037.4]
  wire [31:0] f_13_io_a_bits; // @[TensorAlu.scala 83:36:@22037.4]
  wire  f_13_io_b_valid; // @[TensorAlu.scala 83:36:@22037.4]
  wire [31:0] f_13_io_b_bits; // @[TensorAlu.scala 83:36:@22037.4]
  wire  f_13_io_y_valid; // @[TensorAlu.scala 83:36:@22037.4]
  wire [31:0] f_13_io_y_bits; // @[TensorAlu.scala 83:36:@22037.4]
  wire  f_14_clock; // @[TensorAlu.scala 83:36:@22040.4]
  wire [2:0] f_14_io_opcode; // @[TensorAlu.scala 83:36:@22040.4]
  wire  f_14_io_a_valid; // @[TensorAlu.scala 83:36:@22040.4]
  wire [31:0] f_14_io_a_bits; // @[TensorAlu.scala 83:36:@22040.4]
  wire  f_14_io_b_valid; // @[TensorAlu.scala 83:36:@22040.4]
  wire [31:0] f_14_io_b_bits; // @[TensorAlu.scala 83:36:@22040.4]
  wire  f_14_io_y_valid; // @[TensorAlu.scala 83:36:@22040.4]
  wire [31:0] f_14_io_y_bits; // @[TensorAlu.scala 83:36:@22040.4]
  wire  f_15_clock; // @[TensorAlu.scala 83:36:@22043.4]
  wire [2:0] f_15_io_opcode; // @[TensorAlu.scala 83:36:@22043.4]
  wire  f_15_io_a_valid; // @[TensorAlu.scala 83:36:@22043.4]
  wire [31:0] f_15_io_a_bits; // @[TensorAlu.scala 83:36:@22043.4]
  wire  f_15_io_b_valid; // @[TensorAlu.scala 83:36:@22043.4]
  wire [31:0] f_15_io_b_bits; // @[TensorAlu.scala 83:36:@22043.4]
  wire  f_15_io_y_valid; // @[TensorAlu.scala 83:36:@22043.4]
  wire [31:0] f_15_io_y_bits; // @[TensorAlu.scala 83:36:@22043.4]
  wire  valid_1; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22060.4]
  wire  valid_0; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22052.4]
  wire  valid_3; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22076.4]
  wire  valid_2; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22068.4]
  wire  valid_5; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22092.4]
  wire  valid_4; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22084.4]
  wire  valid_7; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22108.4]
  wire  valid_6; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22100.4]
  wire [7:0] _T_1686; // @[TensorAlu.scala 95:32:@22181.4]
  wire  valid_9; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22124.4]
  wire  valid_8; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22116.4]
  wire  valid_11; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22140.4]
  wire  valid_10; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22132.4]
  wire  valid_13; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22156.4]
  wire  valid_12; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22148.4]
  wire  valid_15; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22172.4]
  wire  valid_14; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22164.4]
  wire [15:0] _T_1694; // @[TensorAlu.scala 95:32:@22189.4]
  wire [15:0] _T_1695; // @[TensorAlu.scala 95:39:@22190.4]
  AluReg f_0 ( // @[TensorAlu.scala 83:36:@21998.4]
    .clock(f_0_clock),
    .io_opcode(f_0_io_opcode),
    .io_a_valid(f_0_io_a_valid),
    .io_a_bits(f_0_io_a_bits),
    .io_b_valid(f_0_io_b_valid),
    .io_b_bits(f_0_io_b_bits),
    .io_y_valid(f_0_io_y_valid),
    .io_y_bits(f_0_io_y_bits)
  );
  AluReg f_1 ( // @[TensorAlu.scala 83:36:@22001.4]
    .clock(f_1_clock),
    .io_opcode(f_1_io_opcode),
    .io_a_valid(f_1_io_a_valid),
    .io_a_bits(f_1_io_a_bits),
    .io_b_valid(f_1_io_b_valid),
    .io_b_bits(f_1_io_b_bits),
    .io_y_valid(f_1_io_y_valid),
    .io_y_bits(f_1_io_y_bits)
  );
  AluReg f_2 ( // @[TensorAlu.scala 83:36:@22004.4]
    .clock(f_2_clock),
    .io_opcode(f_2_io_opcode),
    .io_a_valid(f_2_io_a_valid),
    .io_a_bits(f_2_io_a_bits),
    .io_b_valid(f_2_io_b_valid),
    .io_b_bits(f_2_io_b_bits),
    .io_y_valid(f_2_io_y_valid),
    .io_y_bits(f_2_io_y_bits)
  );
  AluReg f_3 ( // @[TensorAlu.scala 83:36:@22007.4]
    .clock(f_3_clock),
    .io_opcode(f_3_io_opcode),
    .io_a_valid(f_3_io_a_valid),
    .io_a_bits(f_3_io_a_bits),
    .io_b_valid(f_3_io_b_valid),
    .io_b_bits(f_3_io_b_bits),
    .io_y_valid(f_3_io_y_valid),
    .io_y_bits(f_3_io_y_bits)
  );
  AluReg f_4 ( // @[TensorAlu.scala 83:36:@22010.4]
    .clock(f_4_clock),
    .io_opcode(f_4_io_opcode),
    .io_a_valid(f_4_io_a_valid),
    .io_a_bits(f_4_io_a_bits),
    .io_b_valid(f_4_io_b_valid),
    .io_b_bits(f_4_io_b_bits),
    .io_y_valid(f_4_io_y_valid),
    .io_y_bits(f_4_io_y_bits)
  );
  AluReg f_5 ( // @[TensorAlu.scala 83:36:@22013.4]
    .clock(f_5_clock),
    .io_opcode(f_5_io_opcode),
    .io_a_valid(f_5_io_a_valid),
    .io_a_bits(f_5_io_a_bits),
    .io_b_valid(f_5_io_b_valid),
    .io_b_bits(f_5_io_b_bits),
    .io_y_valid(f_5_io_y_valid),
    .io_y_bits(f_5_io_y_bits)
  );
  AluReg f_6 ( // @[TensorAlu.scala 83:36:@22016.4]
    .clock(f_6_clock),
    .io_opcode(f_6_io_opcode),
    .io_a_valid(f_6_io_a_valid),
    .io_a_bits(f_6_io_a_bits),
    .io_b_valid(f_6_io_b_valid),
    .io_b_bits(f_6_io_b_bits),
    .io_y_valid(f_6_io_y_valid),
    .io_y_bits(f_6_io_y_bits)
  );
  AluReg f_7 ( // @[TensorAlu.scala 83:36:@22019.4]
    .clock(f_7_clock),
    .io_opcode(f_7_io_opcode),
    .io_a_valid(f_7_io_a_valid),
    .io_a_bits(f_7_io_a_bits),
    .io_b_valid(f_7_io_b_valid),
    .io_b_bits(f_7_io_b_bits),
    .io_y_valid(f_7_io_y_valid),
    .io_y_bits(f_7_io_y_bits)
  );
  AluReg f_8 ( // @[TensorAlu.scala 83:36:@22022.4]
    .clock(f_8_clock),
    .io_opcode(f_8_io_opcode),
    .io_a_valid(f_8_io_a_valid),
    .io_a_bits(f_8_io_a_bits),
    .io_b_valid(f_8_io_b_valid),
    .io_b_bits(f_8_io_b_bits),
    .io_y_valid(f_8_io_y_valid),
    .io_y_bits(f_8_io_y_bits)
  );
  AluReg f_9 ( // @[TensorAlu.scala 83:36:@22025.4]
    .clock(f_9_clock),
    .io_opcode(f_9_io_opcode),
    .io_a_valid(f_9_io_a_valid),
    .io_a_bits(f_9_io_a_bits),
    .io_b_valid(f_9_io_b_valid),
    .io_b_bits(f_9_io_b_bits),
    .io_y_valid(f_9_io_y_valid),
    .io_y_bits(f_9_io_y_bits)
  );
  AluReg f_10 ( // @[TensorAlu.scala 83:36:@22028.4]
    .clock(f_10_clock),
    .io_opcode(f_10_io_opcode),
    .io_a_valid(f_10_io_a_valid),
    .io_a_bits(f_10_io_a_bits),
    .io_b_valid(f_10_io_b_valid),
    .io_b_bits(f_10_io_b_bits),
    .io_y_valid(f_10_io_y_valid),
    .io_y_bits(f_10_io_y_bits)
  );
  AluReg f_11 ( // @[TensorAlu.scala 83:36:@22031.4]
    .clock(f_11_clock),
    .io_opcode(f_11_io_opcode),
    .io_a_valid(f_11_io_a_valid),
    .io_a_bits(f_11_io_a_bits),
    .io_b_valid(f_11_io_b_valid),
    .io_b_bits(f_11_io_b_bits),
    .io_y_valid(f_11_io_y_valid),
    .io_y_bits(f_11_io_y_bits)
  );
  AluReg f_12 ( // @[TensorAlu.scala 83:36:@22034.4]
    .clock(f_12_clock),
    .io_opcode(f_12_io_opcode),
    .io_a_valid(f_12_io_a_valid),
    .io_a_bits(f_12_io_a_bits),
    .io_b_valid(f_12_io_b_valid),
    .io_b_bits(f_12_io_b_bits),
    .io_y_valid(f_12_io_y_valid),
    .io_y_bits(f_12_io_y_bits)
  );
  AluReg f_13 ( // @[TensorAlu.scala 83:36:@22037.4]
    .clock(f_13_clock),
    .io_opcode(f_13_io_opcode),
    .io_a_valid(f_13_io_a_valid),
    .io_a_bits(f_13_io_a_bits),
    .io_b_valid(f_13_io_b_valid),
    .io_b_bits(f_13_io_b_bits),
    .io_y_valid(f_13_io_y_valid),
    .io_y_bits(f_13_io_y_bits)
  );
  AluReg f_14 ( // @[TensorAlu.scala 83:36:@22040.4]
    .clock(f_14_clock),
    .io_opcode(f_14_io_opcode),
    .io_a_valid(f_14_io_a_valid),
    .io_a_bits(f_14_io_a_bits),
    .io_b_valid(f_14_io_b_valid),
    .io_b_bits(f_14_io_b_bits),
    .io_y_valid(f_14_io_y_valid),
    .io_y_bits(f_14_io_y_bits)
  );
  AluReg f_15 ( // @[TensorAlu.scala 83:36:@22043.4]
    .clock(f_15_clock),
    .io_opcode(f_15_io_opcode),
    .io_a_valid(f_15_io_a_valid),
    .io_a_bits(f_15_io_a_bits),
    .io_b_valid(f_15_io_b_valid),
    .io_b_bits(f_15_io_b_bits),
    .io_y_valid(f_15_io_y_valid),
    .io_y_bits(f_15_io_y_bits)
  );
  assign valid_1 = f_1_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22060.4]
  assign valid_0 = f_0_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22052.4]
  assign valid_3 = f_3_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22076.4]
  assign valid_2 = f_2_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22068.4]
  assign valid_5 = f_5_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22092.4]
  assign valid_4 = f_4_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22084.4]
  assign valid_7 = f_7_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22108.4]
  assign valid_6 = f_6_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22100.4]
  assign _T_1686 = {valid_7,valid_6,valid_5,valid_4,valid_3,valid_2,valid_1,valid_0}; // @[TensorAlu.scala 95:32:@22181.4]
  assign valid_9 = f_9_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22124.4]
  assign valid_8 = f_8_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22116.4]
  assign valid_11 = f_11_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22140.4]
  assign valid_10 = f_10_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22132.4]
  assign valid_13 = f_13_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22156.4]
  assign valid_12 = f_12_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22148.4]
  assign valid_15 = f_15_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22172.4]
  assign valid_14 = f_14_io_y_valid; // @[TensorAlu.scala 84:19:@22046.4 TensorAlu.scala 91:14:@22164.4]
  assign _T_1694 = {valid_15,valid_14,valid_13,valid_12,valid_11,valid_10,valid_9,valid_8,_T_1686}; // @[TensorAlu.scala 95:32:@22189.4]
  assign _T_1695 = ~ _T_1694; // @[TensorAlu.scala 95:39:@22190.4]
  assign io_acc_y_data_valid = _T_1695 == 16'h0; // @[TensorAlu.scala 95:23:@22192.4]
  assign io_acc_y_data_bits_0_0 = f_0_io_y_bits; // @[TensorAlu.scala 92:30:@22053.4]
  assign io_acc_y_data_bits_0_1 = f_1_io_y_bits; // @[TensorAlu.scala 92:30:@22061.4]
  assign io_acc_y_data_bits_0_2 = f_2_io_y_bits; // @[TensorAlu.scala 92:30:@22069.4]
  assign io_acc_y_data_bits_0_3 = f_3_io_y_bits; // @[TensorAlu.scala 92:30:@22077.4]
  assign io_acc_y_data_bits_0_4 = f_4_io_y_bits; // @[TensorAlu.scala 92:30:@22085.4]
  assign io_acc_y_data_bits_0_5 = f_5_io_y_bits; // @[TensorAlu.scala 92:30:@22093.4]
  assign io_acc_y_data_bits_0_6 = f_6_io_y_bits; // @[TensorAlu.scala 92:30:@22101.4]
  assign io_acc_y_data_bits_0_7 = f_7_io_y_bits; // @[TensorAlu.scala 92:30:@22109.4]
  assign io_acc_y_data_bits_0_8 = f_8_io_y_bits; // @[TensorAlu.scala 92:30:@22117.4]
  assign io_acc_y_data_bits_0_9 = f_9_io_y_bits; // @[TensorAlu.scala 92:30:@22125.4]
  assign io_acc_y_data_bits_0_10 = f_10_io_y_bits; // @[TensorAlu.scala 92:30:@22133.4]
  assign io_acc_y_data_bits_0_11 = f_11_io_y_bits; // @[TensorAlu.scala 92:30:@22141.4]
  assign io_acc_y_data_bits_0_12 = f_12_io_y_bits; // @[TensorAlu.scala 92:30:@22149.4]
  assign io_acc_y_data_bits_0_13 = f_13_io_y_bits; // @[TensorAlu.scala 92:30:@22157.4]
  assign io_acc_y_data_bits_0_14 = f_14_io_y_bits; // @[TensorAlu.scala 92:30:@22165.4]
  assign io_acc_y_data_bits_0_15 = f_15_io_y_bits; // @[TensorAlu.scala 92:30:@22173.4]
  assign io_out_data_valid = _T_1695 == 16'h0; // @[TensorAlu.scala 96:21:@22210.4]
  assign io_out_data_bits_0_0 = f_0_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22054.4]
  assign io_out_data_bits_0_1 = f_1_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22062.4]
  assign io_out_data_bits_0_2 = f_2_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22070.4]
  assign io_out_data_bits_0_3 = f_3_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22078.4]
  assign io_out_data_bits_0_4 = f_4_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22086.4]
  assign io_out_data_bits_0_5 = f_5_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22094.4]
  assign io_out_data_bits_0_6 = f_6_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22102.4]
  assign io_out_data_bits_0_7 = f_7_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22110.4]
  assign io_out_data_bits_0_8 = f_8_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22118.4]
  assign io_out_data_bits_0_9 = f_9_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22126.4]
  assign io_out_data_bits_0_10 = f_10_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22134.4]
  assign io_out_data_bits_0_11 = f_11_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22142.4]
  assign io_out_data_bits_0_12 = f_12_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22150.4]
  assign io_out_data_bits_0_13 = f_13_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22158.4]
  assign io_out_data_bits_0_14 = f_14_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22166.4]
  assign io_out_data_bits_0_15 = f_15_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22174.4]
  assign f_0_clock = clock; // @[:@21999.4]
  assign f_0_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22047.4]
  assign f_0_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22048.4]
  assign f_0_io_a_bits = io_acc_a_data_bits_0_0; // @[TensorAlu.scala 88:20:@22049.4]
  assign f_0_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22050.4]
  assign f_0_io_b_bits = io_acc_b_data_bits_0_0; // @[TensorAlu.scala 90:20:@22051.4]
  assign f_1_clock = clock; // @[:@22002.4]
  assign f_1_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22055.4]
  assign f_1_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22056.4]
  assign f_1_io_a_bits = io_acc_a_data_bits_0_1; // @[TensorAlu.scala 88:20:@22057.4]
  assign f_1_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22058.4]
  assign f_1_io_b_bits = io_acc_b_data_bits_0_1; // @[TensorAlu.scala 90:20:@22059.4]
  assign f_2_clock = clock; // @[:@22005.4]
  assign f_2_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22063.4]
  assign f_2_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22064.4]
  assign f_2_io_a_bits = io_acc_a_data_bits_0_2; // @[TensorAlu.scala 88:20:@22065.4]
  assign f_2_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22066.4]
  assign f_2_io_b_bits = io_acc_b_data_bits_0_2; // @[TensorAlu.scala 90:20:@22067.4]
  assign f_3_clock = clock; // @[:@22008.4]
  assign f_3_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22071.4]
  assign f_3_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22072.4]
  assign f_3_io_a_bits = io_acc_a_data_bits_0_3; // @[TensorAlu.scala 88:20:@22073.4]
  assign f_3_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22074.4]
  assign f_3_io_b_bits = io_acc_b_data_bits_0_3; // @[TensorAlu.scala 90:20:@22075.4]
  assign f_4_clock = clock; // @[:@22011.4]
  assign f_4_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22079.4]
  assign f_4_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22080.4]
  assign f_4_io_a_bits = io_acc_a_data_bits_0_4; // @[TensorAlu.scala 88:20:@22081.4]
  assign f_4_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22082.4]
  assign f_4_io_b_bits = io_acc_b_data_bits_0_4; // @[TensorAlu.scala 90:20:@22083.4]
  assign f_5_clock = clock; // @[:@22014.4]
  assign f_5_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22087.4]
  assign f_5_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22088.4]
  assign f_5_io_a_bits = io_acc_a_data_bits_0_5; // @[TensorAlu.scala 88:20:@22089.4]
  assign f_5_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22090.4]
  assign f_5_io_b_bits = io_acc_b_data_bits_0_5; // @[TensorAlu.scala 90:20:@22091.4]
  assign f_6_clock = clock; // @[:@22017.4]
  assign f_6_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22095.4]
  assign f_6_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22096.4]
  assign f_6_io_a_bits = io_acc_a_data_bits_0_6; // @[TensorAlu.scala 88:20:@22097.4]
  assign f_6_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22098.4]
  assign f_6_io_b_bits = io_acc_b_data_bits_0_6; // @[TensorAlu.scala 90:20:@22099.4]
  assign f_7_clock = clock; // @[:@22020.4]
  assign f_7_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22103.4]
  assign f_7_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22104.4]
  assign f_7_io_a_bits = io_acc_a_data_bits_0_7; // @[TensorAlu.scala 88:20:@22105.4]
  assign f_7_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22106.4]
  assign f_7_io_b_bits = io_acc_b_data_bits_0_7; // @[TensorAlu.scala 90:20:@22107.4]
  assign f_8_clock = clock; // @[:@22023.4]
  assign f_8_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22111.4]
  assign f_8_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22112.4]
  assign f_8_io_a_bits = io_acc_a_data_bits_0_8; // @[TensorAlu.scala 88:20:@22113.4]
  assign f_8_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22114.4]
  assign f_8_io_b_bits = io_acc_b_data_bits_0_8; // @[TensorAlu.scala 90:20:@22115.4]
  assign f_9_clock = clock; // @[:@22026.4]
  assign f_9_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22119.4]
  assign f_9_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22120.4]
  assign f_9_io_a_bits = io_acc_a_data_bits_0_9; // @[TensorAlu.scala 88:20:@22121.4]
  assign f_9_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22122.4]
  assign f_9_io_b_bits = io_acc_b_data_bits_0_9; // @[TensorAlu.scala 90:20:@22123.4]
  assign f_10_clock = clock; // @[:@22029.4]
  assign f_10_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22127.4]
  assign f_10_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22128.4]
  assign f_10_io_a_bits = io_acc_a_data_bits_0_10; // @[TensorAlu.scala 88:20:@22129.4]
  assign f_10_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22130.4]
  assign f_10_io_b_bits = io_acc_b_data_bits_0_10; // @[TensorAlu.scala 90:20:@22131.4]
  assign f_11_clock = clock; // @[:@22032.4]
  assign f_11_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22135.4]
  assign f_11_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22136.4]
  assign f_11_io_a_bits = io_acc_a_data_bits_0_11; // @[TensorAlu.scala 88:20:@22137.4]
  assign f_11_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22138.4]
  assign f_11_io_b_bits = io_acc_b_data_bits_0_11; // @[TensorAlu.scala 90:20:@22139.4]
  assign f_12_clock = clock; // @[:@22035.4]
  assign f_12_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22143.4]
  assign f_12_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22144.4]
  assign f_12_io_a_bits = io_acc_a_data_bits_0_12; // @[TensorAlu.scala 88:20:@22145.4]
  assign f_12_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22146.4]
  assign f_12_io_b_bits = io_acc_b_data_bits_0_12; // @[TensorAlu.scala 90:20:@22147.4]
  assign f_13_clock = clock; // @[:@22038.4]
  assign f_13_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22151.4]
  assign f_13_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22152.4]
  assign f_13_io_a_bits = io_acc_a_data_bits_0_13; // @[TensorAlu.scala 88:20:@22153.4]
  assign f_13_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22154.4]
  assign f_13_io_b_bits = io_acc_b_data_bits_0_13; // @[TensorAlu.scala 90:20:@22155.4]
  assign f_14_clock = clock; // @[:@22041.4]
  assign f_14_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22159.4]
  assign f_14_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22160.4]
  assign f_14_io_a_bits = io_acc_a_data_bits_0_14; // @[TensorAlu.scala 88:20:@22161.4]
  assign f_14_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22162.4]
  assign f_14_io_b_bits = io_acc_b_data_bits_0_14; // @[TensorAlu.scala 90:20:@22163.4]
  assign f_15_clock = clock; // @[:@22044.4]
  assign f_15_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22167.4]
  assign f_15_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22168.4]
  assign f_15_io_a_bits = io_acc_a_data_bits_0_15; // @[TensorAlu.scala 88:20:@22169.4]
  assign f_15_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22170.4]
  assign f_15_io_b_bits = io_acc_b_data_bits_0_15; // @[TensorAlu.scala 90:20:@22171.4]
endmodule
module TensorAlu( // @[:@22212.2]
  input          clock, // @[:@22213.4]
  input          reset, // @[:@22214.4]
  input          io_start, // @[:@22215.4]
  output         io_done, // @[:@22215.4]
  input  [127:0] io_inst, // @[:@22215.4]
  output         io_uop_idx_valid, // @[:@22215.4]
  output [10:0]  io_uop_idx_bits, // @[:@22215.4]
  input          io_uop_data_valid, // @[:@22215.4]
  input  [10:0]  io_uop_data_bits_u1, // @[:@22215.4]
  input  [10:0]  io_uop_data_bits_u0, // @[:@22215.4]
  output         io_acc_rd_idx_valid, // @[:@22215.4]
  output [10:0]  io_acc_rd_idx_bits, // @[:@22215.4]
  input          io_acc_rd_data_valid, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_0, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_1, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_2, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_3, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_4, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_5, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_6, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_7, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_8, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_9, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_10, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_11, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_12, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_13, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_14, // @[:@22215.4]
  input  [31:0]  io_acc_rd_data_bits_0_15, // @[:@22215.4]
  output         io_acc_wr_valid, // @[:@22215.4]
  output [10:0]  io_acc_wr_bits_idx, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_0, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_1, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_2, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_3, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_4, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_5, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_6, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_7, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_8, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_9, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_10, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_11, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_12, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_13, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_14, // @[:@22215.4]
  output [31:0]  io_acc_wr_bits_data_0_15, // @[:@22215.4]
  output         io_out_wr_valid, // @[:@22215.4]
  output [10:0]  io_out_wr_bits_idx, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_0, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_1, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_2, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_3, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_4, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_5, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_6, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_7, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_8, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_9, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_10, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_11, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_12, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_13, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_14, // @[:@22215.4]
  output [7:0]   io_out_wr_bits_data_0_15 // @[:@22215.4]
);
  wire  alu_clock; // @[TensorAlu.scala 119:19:@22218.4]
  wire [2:0] alu_io_opcode; // @[TensorAlu.scala 119:19:@22218.4]
  wire  alu_io_acc_a_data_valid; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_0; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_1; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_2; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_3; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_4; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_5; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_6; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_7; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_8; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_9; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_10; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_11; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_12; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_13; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_14; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_a_data_bits_0_15; // @[TensorAlu.scala 119:19:@22218.4]
  wire  alu_io_acc_b_data_valid; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_0; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_1; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_2; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_3; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_4; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_5; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_6; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_7; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_8; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_9; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_10; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_11; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_12; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_13; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_14; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_b_data_bits_0_15; // @[TensorAlu.scala 119:19:@22218.4]
  wire  alu_io_acc_y_data_valid; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_0; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_1; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_2; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_3; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_4; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_5; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_6; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_7; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_8; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_9; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_10; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_11; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_12; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_13; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_14; // @[TensorAlu.scala 119:19:@22218.4]
  wire [31:0] alu_io_acc_y_data_bits_0_15; // @[TensorAlu.scala 119:19:@22218.4]
  wire  alu_io_out_data_valid; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_0; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_1; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_2; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_3; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_4; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_5; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_6; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_7; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_8; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_9; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_10; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_11; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_12; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_13; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_14; // @[TensorAlu.scala 119:19:@22218.4]
  wire [7:0] alu_io_out_data_bits_0_15; // @[TensorAlu.scala 119:19:@22218.4]
  reg [2:0] state; // @[TensorAlu.scala 118:22:@22217.4]
  reg [31:0] _RAND_0;
  wire [12:0] dec_uop_begin; // @[TensorAlu.scala 120:29:@22236.4]
  wire [13:0] dec_uop_end; // @[TensorAlu.scala 120:29:@22238.4]
  wire [13:0] dec_lp_0; // @[TensorAlu.scala 120:29:@22240.4]
  wire [13:0] dec_lp_1; // @[TensorAlu.scala 120:29:@22242.4]
  wire [10:0] dec_dst_0; // @[TensorAlu.scala 120:29:@22246.4]
  wire [10:0] dec_dst_1; // @[TensorAlu.scala 120:29:@22248.4]
  wire [10:0] dec_src_0; // @[TensorAlu.scala 120:29:@22250.4]
  wire [10:0] dec_src_1; // @[TensorAlu.scala 120:29:@22252.4]
  wire [1:0] dec_alu_op; // @[TensorAlu.scala 120:29:@22254.4]
  wire  dec_alu_use_imm; // @[TensorAlu.scala 120:29:@22256.4]
  wire [15:0] dec_alu_imm; // @[TensorAlu.scala 120:29:@22258.4]
  reg [13:0] uop_idx; // @[TensorAlu.scala 121:20:@22262.4]
  reg [31:0] _RAND_1;
  reg [13:0] uop_dst; // @[TensorAlu.scala 123:20:@22263.4]
  reg [31:0] _RAND_2;
  reg [13:0] uop_src; // @[TensorAlu.scala 124:20:@22264.4]
  reg [31:0] _RAND_3;
  reg [13:0] cnt_o; // @[TensorAlu.scala 125:18:@22265.4]
  reg [31:0] _RAND_4;
  reg [13:0] dst_o; // @[TensorAlu.scala 126:18:@22266.4]
  reg [31:0] _RAND_5;
  reg [13:0] src_o; // @[TensorAlu.scala 127:18:@22267.4]
  reg [31:0] _RAND_6;
  reg [13:0] cnt_i; // @[TensorAlu.scala 128:18:@22268.4]
  reg [31:0] _RAND_7;
  reg [13:0] dst_i; // @[TensorAlu.scala 129:18:@22269.4]
  reg [31:0] _RAND_8;
  reg [13:0] src_i; // @[TensorAlu.scala 130:18:@22270.4]
  reg [31:0] _RAND_9;
  wire  _T_1440; // @[TensorAlu.scala 132:11:@22271.4]
  wire  _T_1441; // @[TensorAlu.scala 132:20:@22272.4]
  wire [14:0] _T_1443; // @[TensorAlu.scala 134:27:@22273.4]
  wire [14:0] _T_1444; // @[TensorAlu.scala 134:27:@22274.4]
  wire [13:0] _T_1445; // @[TensorAlu.scala 134:27:@22275.4]
  wire  _T_1446; // @[TensorAlu.scala 134:14:@22276.4]
  wire  _T_1447; // @[TensorAlu.scala 133:29:@22277.4]
  wire [14:0] _T_1449; // @[TensorAlu.scala 135:27:@22278.4]
  wire [14:0] _T_1450; // @[TensorAlu.scala 135:27:@22279.4]
  wire [13:0] _T_1451; // @[TensorAlu.scala 135:27:@22280.4]
  wire  _T_1452; // @[TensorAlu.scala 135:14:@22281.4]
  wire  _T_1453; // @[TensorAlu.scala 134:34:@22282.4]
  wire [14:0] _T_1455; // @[TensorAlu.scala 136:28:@22283.4]
  wire [14:0] _T_1456; // @[TensorAlu.scala 136:28:@22284.4]
  wire [13:0] _T_1457; // @[TensorAlu.scala 136:28:@22285.4]
  wire  _T_1458; // @[TensorAlu.scala 136:16:@22286.4]
  wire  _T_1459; // @[Conditional.scala 37:30:@22288.4]
  wire [2:0] _GEN_0; // @[TensorAlu.scala 140:22:@22290.6]
  wire  _T_1460; // @[Conditional.scala 37:30:@22295.6]
  wire  _T_1461; // @[Conditional.scala 37:30:@22300.8]
  wire  _T_1462; // @[Conditional.scala 37:30:@22305.10]
  wire  _T_1463; // @[Conditional.scala 37:30:@22310.12]
  wire  _T_1464; // @[Conditional.scala 37:30:@22315.14]
  wire  _T_1475; // @[TensorAlu.scala 159:38:@22326.18]
  wire  _T_1481; // @[TensorAlu.scala 160:40:@22331.18]
  wire [2:0] _GEN_1; // @[TensorAlu.scala 161:42:@22332.18]
  wire [2:0] _GEN_2; // @[TensorAlu.scala 157:35:@22317.16]
  wire [2:0] _GEN_3; // @[Conditional.scala 39:67:@22316.14]
  wire [2:0] _GEN_4; // @[Conditional.scala 39:67:@22311.12]
  wire [2:0] _GEN_5; // @[Conditional.scala 39:67:@22306.10]
  wire [2:0] _GEN_6; // @[Conditional.scala 39:67:@22301.8]
  wire [2:0] _GEN_7; // @[Conditional.scala 39:67:@22296.6]
  wire [2:0] _GEN_8; // @[Conditional.scala 40:58:@22289.4]
  wire  _T_1482; // @[TensorAlu.scala 171:11:@22340.4]
  wire  _T_1490; // @[TensorAlu.scala 173:31:@22347.4]
  wire  _T_1491; // @[TensorAlu.scala 171:21:@22348.4]
  wire [14:0] _T_1495; // @[TensorAlu.scala 177:24:@22356.8]
  wire [13:0] _T_1496; // @[TensorAlu.scala 177:24:@22357.8]
  wire [13:0] _GEN_9; // @[TensorAlu.scala 176:55:@22355.6]
  wire  _T_1514; // @[TensorAlu.scala 187:33:@22378.6]
  wire [14:0] _T_1516; // @[TensorAlu.scala 189:20:@22380.8]
  wire [13:0] _T_1517; // @[TensorAlu.scala 189:20:@22381.8]
  wire [13:0] _GEN_28; // @[TensorAlu.scala 190:20:@22383.8]
  wire [14:0] _T_1518; // @[TensorAlu.scala 190:20:@22383.8]
  wire [13:0] _T_1519; // @[TensorAlu.scala 190:20:@22384.8]
  wire [13:0] _GEN_29; // @[TensorAlu.scala 191:20:@22386.8]
  wire [14:0] _T_1520; // @[TensorAlu.scala 191:20:@22386.8]
  wire [13:0] _T_1521; // @[TensorAlu.scala 191:20:@22387.8]
  wire [13:0] _GEN_11; // @[TensorAlu.scala 188:33:@22379.6]
  wire [13:0] _GEN_12; // @[TensorAlu.scala 188:33:@22379.6]
  wire [13:0] _GEN_13; // @[TensorAlu.scala 188:33:@22379.6]
  wire  _T_1526; // @[TensorAlu.scala 198:20:@22397.6]
  wire  _T_1527; // @[TensorAlu.scala 198:42:@22398.6]
  wire  _T_1528; // @[TensorAlu.scala 198:33:@22399.6]
  wire [14:0] _T_1539; // @[TensorAlu.scala 203:20:@22414.10]
  wire [13:0] _T_1540; // @[TensorAlu.scala 203:20:@22415.10]
  wire [13:0] _GEN_30; // @[TensorAlu.scala 204:20:@22417.10]
  wire [14:0] _T_1541; // @[TensorAlu.scala 204:20:@22417.10]
  wire [13:0] _T_1542; // @[TensorAlu.scala 204:20:@22418.10]
  wire [13:0] _GEN_31; // @[TensorAlu.scala 205:20:@22420.10]
  wire [14:0] _T_1543; // @[TensorAlu.scala 205:20:@22420.10]
  wire [13:0] _T_1544; // @[TensorAlu.scala 205:20:@22421.10]
  wire [13:0] _GEN_17; // @[TensorAlu.scala 202:84:@22413.8]
  wire [13:0] _GEN_18; // @[TensorAlu.scala 202:84:@22413.8]
  wire [13:0] _GEN_19; // @[TensorAlu.scala 202:84:@22413.8]
  wire [13:0] _GEN_20; // @[TensorAlu.scala 198:56:@22400.6]
  wire [13:0] _GEN_21; // @[TensorAlu.scala 198:56:@22400.6]
  wire [13:0] _GEN_22; // @[TensorAlu.scala 198:56:@22400.6]
  wire  _T_1545; // @[TensorAlu.scala 208:14:@22424.4]
  wire  _T_1546; // @[TensorAlu.scala 208:30:@22425.4]
  wire [13:0] _GEN_32; // @[TensorAlu.scala 209:36:@22427.6]
  wire [14:0] _T_1547; // @[TensorAlu.scala 209:36:@22427.6]
  wire [13:0] _T_1548; // @[TensorAlu.scala 209:36:@22428.6]
  wire [13:0] _GEN_33; // @[TensorAlu.scala 210:36:@22430.6]
  wire [14:0] _T_1549; // @[TensorAlu.scala 210:36:@22430.6]
  wire [13:0] _T_1550; // @[TensorAlu.scala 210:36:@22431.6]
  wire  _T_1552; // @[TensorAlu.scala 218:32:@22437.4]
  wire  _T_1553; // @[TensorAlu.scala 218:58:@22438.4]
  wire  _T_1554; // @[TensorAlu.scala 218:77:@22439.4]
  wire  _T_1555; // @[TensorAlu.scala 218:75:@22440.4]
  wire [13:0] _T_1558; // @[TensorAlu.scala 219:28:@22444.4]
  wire  _T_1863; // @[TensorAlu.scala 226:27:@22449.4]
  wire [31:0] _T_1866; // @[Cat.scala 30:58:@22451.4]
  wire [31:0] tensorImm_data_bits_0_0; // @[TensorAlu.scala 226:15:@22452.4]
  wire [2:0] _GEN_34; // @[TensorAlu.scala 232:26:@22529.4]
  wire  isSHR; // @[TensorAlu.scala 232:26:@22529.4]
  wire  neg_shift; // @[TensorAlu.scala 233:25:@22531.4]
  wire [1:0] _T_1945; // @[TensorAlu.scala 234:40:@22532.4]
  wire  _T_1949; // @[TensorAlu.scala 240:26:@22555.4]
  AluVector alu ( // @[TensorAlu.scala 119:19:@22218.4]
    .clock(alu_clock),
    .io_opcode(alu_io_opcode),
    .io_acc_a_data_valid(alu_io_acc_a_data_valid),
    .io_acc_a_data_bits_0_0(alu_io_acc_a_data_bits_0_0),
    .io_acc_a_data_bits_0_1(alu_io_acc_a_data_bits_0_1),
    .io_acc_a_data_bits_0_2(alu_io_acc_a_data_bits_0_2),
    .io_acc_a_data_bits_0_3(alu_io_acc_a_data_bits_0_3),
    .io_acc_a_data_bits_0_4(alu_io_acc_a_data_bits_0_4),
    .io_acc_a_data_bits_0_5(alu_io_acc_a_data_bits_0_5),
    .io_acc_a_data_bits_0_6(alu_io_acc_a_data_bits_0_6),
    .io_acc_a_data_bits_0_7(alu_io_acc_a_data_bits_0_7),
    .io_acc_a_data_bits_0_8(alu_io_acc_a_data_bits_0_8),
    .io_acc_a_data_bits_0_9(alu_io_acc_a_data_bits_0_9),
    .io_acc_a_data_bits_0_10(alu_io_acc_a_data_bits_0_10),
    .io_acc_a_data_bits_0_11(alu_io_acc_a_data_bits_0_11),
    .io_acc_a_data_bits_0_12(alu_io_acc_a_data_bits_0_12),
    .io_acc_a_data_bits_0_13(alu_io_acc_a_data_bits_0_13),
    .io_acc_a_data_bits_0_14(alu_io_acc_a_data_bits_0_14),
    .io_acc_a_data_bits_0_15(alu_io_acc_a_data_bits_0_15),
    .io_acc_b_data_valid(alu_io_acc_b_data_valid),
    .io_acc_b_data_bits_0_0(alu_io_acc_b_data_bits_0_0),
    .io_acc_b_data_bits_0_1(alu_io_acc_b_data_bits_0_1),
    .io_acc_b_data_bits_0_2(alu_io_acc_b_data_bits_0_2),
    .io_acc_b_data_bits_0_3(alu_io_acc_b_data_bits_0_3),
    .io_acc_b_data_bits_0_4(alu_io_acc_b_data_bits_0_4),
    .io_acc_b_data_bits_0_5(alu_io_acc_b_data_bits_0_5),
    .io_acc_b_data_bits_0_6(alu_io_acc_b_data_bits_0_6),
    .io_acc_b_data_bits_0_7(alu_io_acc_b_data_bits_0_7),
    .io_acc_b_data_bits_0_8(alu_io_acc_b_data_bits_0_8),
    .io_acc_b_data_bits_0_9(alu_io_acc_b_data_bits_0_9),
    .io_acc_b_data_bits_0_10(alu_io_acc_b_data_bits_0_10),
    .io_acc_b_data_bits_0_11(alu_io_acc_b_data_bits_0_11),
    .io_acc_b_data_bits_0_12(alu_io_acc_b_data_bits_0_12),
    .io_acc_b_data_bits_0_13(alu_io_acc_b_data_bits_0_13),
    .io_acc_b_data_bits_0_14(alu_io_acc_b_data_bits_0_14),
    .io_acc_b_data_bits_0_15(alu_io_acc_b_data_bits_0_15),
    .io_acc_y_data_valid(alu_io_acc_y_data_valid),
    .io_acc_y_data_bits_0_0(alu_io_acc_y_data_bits_0_0),
    .io_acc_y_data_bits_0_1(alu_io_acc_y_data_bits_0_1),
    .io_acc_y_data_bits_0_2(alu_io_acc_y_data_bits_0_2),
    .io_acc_y_data_bits_0_3(alu_io_acc_y_data_bits_0_3),
    .io_acc_y_data_bits_0_4(alu_io_acc_y_data_bits_0_4),
    .io_acc_y_data_bits_0_5(alu_io_acc_y_data_bits_0_5),
    .io_acc_y_data_bits_0_6(alu_io_acc_y_data_bits_0_6),
    .io_acc_y_data_bits_0_7(alu_io_acc_y_data_bits_0_7),
    .io_acc_y_data_bits_0_8(alu_io_acc_y_data_bits_0_8),
    .io_acc_y_data_bits_0_9(alu_io_acc_y_data_bits_0_9),
    .io_acc_y_data_bits_0_10(alu_io_acc_y_data_bits_0_10),
    .io_acc_y_data_bits_0_11(alu_io_acc_y_data_bits_0_11),
    .io_acc_y_data_bits_0_12(alu_io_acc_y_data_bits_0_12),
    .io_acc_y_data_bits_0_13(alu_io_acc_y_data_bits_0_13),
    .io_acc_y_data_bits_0_14(alu_io_acc_y_data_bits_0_14),
    .io_acc_y_data_bits_0_15(alu_io_acc_y_data_bits_0_15),
    .io_out_data_valid(alu_io_out_data_valid),
    .io_out_data_bits_0_0(alu_io_out_data_bits_0_0),
    .io_out_data_bits_0_1(alu_io_out_data_bits_0_1),
    .io_out_data_bits_0_2(alu_io_out_data_bits_0_2),
    .io_out_data_bits_0_3(alu_io_out_data_bits_0_3),
    .io_out_data_bits_0_4(alu_io_out_data_bits_0_4),
    .io_out_data_bits_0_5(alu_io_out_data_bits_0_5),
    .io_out_data_bits_0_6(alu_io_out_data_bits_0_6),
    .io_out_data_bits_0_7(alu_io_out_data_bits_0_7),
    .io_out_data_bits_0_8(alu_io_out_data_bits_0_8),
    .io_out_data_bits_0_9(alu_io_out_data_bits_0_9),
    .io_out_data_bits_0_10(alu_io_out_data_bits_0_10),
    .io_out_data_bits_0_11(alu_io_out_data_bits_0_11),
    .io_out_data_bits_0_12(alu_io_out_data_bits_0_12),
    .io_out_data_bits_0_13(alu_io_out_data_bits_0_13),
    .io_out_data_bits_0_14(alu_io_out_data_bits_0_14),
    .io_out_data_bits_0_15(alu_io_out_data_bits_0_15)
  );
  assign dec_uop_begin = io_inst[20:8]; // @[TensorAlu.scala 120:29:@22236.4]
  assign dec_uop_end = io_inst[34:21]; // @[TensorAlu.scala 120:29:@22238.4]
  assign dec_lp_0 = io_inst[48:35]; // @[TensorAlu.scala 120:29:@22240.4]
  assign dec_lp_1 = io_inst[62:49]; // @[TensorAlu.scala 120:29:@22242.4]
  assign dec_dst_0 = io_inst[74:64]; // @[TensorAlu.scala 120:29:@22246.4]
  assign dec_dst_1 = io_inst[85:75]; // @[TensorAlu.scala 120:29:@22248.4]
  assign dec_src_0 = io_inst[96:86]; // @[TensorAlu.scala 120:29:@22250.4]
  assign dec_src_1 = io_inst[107:97]; // @[TensorAlu.scala 120:29:@22252.4]
  assign dec_alu_op = io_inst[109:108]; // @[TensorAlu.scala 120:29:@22254.4]
  assign dec_alu_use_imm = io_inst[110]; // @[TensorAlu.scala 120:29:@22256.4]
  assign dec_alu_imm = io_inst[126:111]; // @[TensorAlu.scala 120:29:@22258.4]
  assign _T_1440 = state == 3'h5; // @[TensorAlu.scala 132:11:@22271.4]
  assign _T_1441 = _T_1440 & alu_io_out_data_valid; // @[TensorAlu.scala 132:20:@22272.4]
  assign _T_1443 = dec_lp_0 - 14'h1; // @[TensorAlu.scala 134:27:@22273.4]
  assign _T_1444 = $unsigned(_T_1443); // @[TensorAlu.scala 134:27:@22274.4]
  assign _T_1445 = _T_1444[13:0]; // @[TensorAlu.scala 134:27:@22275.4]
  assign _T_1446 = cnt_o == _T_1445; // @[TensorAlu.scala 134:14:@22276.4]
  assign _T_1447 = _T_1441 & _T_1446; // @[TensorAlu.scala 133:29:@22277.4]
  assign _T_1449 = dec_lp_1 - 14'h1; // @[TensorAlu.scala 135:27:@22278.4]
  assign _T_1450 = $unsigned(_T_1449); // @[TensorAlu.scala 135:27:@22279.4]
  assign _T_1451 = _T_1450[13:0]; // @[TensorAlu.scala 135:27:@22280.4]
  assign _T_1452 = cnt_i == _T_1451; // @[TensorAlu.scala 135:14:@22281.4]
  assign _T_1453 = _T_1447 & _T_1452; // @[TensorAlu.scala 134:34:@22282.4]
  assign _T_1455 = dec_uop_end - 14'h1; // @[TensorAlu.scala 136:28:@22283.4]
  assign _T_1456 = $unsigned(_T_1455); // @[TensorAlu.scala 136:28:@22284.4]
  assign _T_1457 = _T_1456[13:0]; // @[TensorAlu.scala 136:28:@22285.4]
  assign _T_1458 = uop_idx == _T_1457; // @[TensorAlu.scala 136:16:@22286.4]
  assign _T_1459 = 3'h0 == state; // @[Conditional.scala 37:30:@22288.4]
  assign _GEN_0 = io_start ? 3'h1 : state; // @[TensorAlu.scala 140:22:@22290.6]
  assign _T_1460 = 3'h1 == state; // @[Conditional.scala 37:30:@22295.6]
  assign _T_1461 = 3'h2 == state; // @[Conditional.scala 37:30:@22300.8]
  assign _T_1462 = 3'h3 == state; // @[Conditional.scala 37:30:@22305.10]
  assign _T_1463 = 3'h4 == state; // @[Conditional.scala 37:30:@22310.12]
  assign _T_1464 = 3'h5 == state; // @[Conditional.scala 37:30:@22315.14]
  assign _T_1475 = _T_1446 & _T_1452; // @[TensorAlu.scala 159:38:@22326.18]
  assign _T_1481 = _T_1475 & _T_1458; // @[TensorAlu.scala 160:40:@22331.18]
  assign _GEN_1 = _T_1481 ? 3'h0 : 3'h1; // @[TensorAlu.scala 161:42:@22332.18]
  assign _GEN_2 = alu_io_out_data_valid ? _GEN_1 : state; // @[TensorAlu.scala 157:35:@22317.16]
  assign _GEN_3 = _T_1464 ? _GEN_2 : state; // @[Conditional.scala 39:67:@22316.14]
  assign _GEN_4 = _T_1463 ? 3'h5 : _GEN_3; // @[Conditional.scala 39:67:@22311.12]
  assign _GEN_5 = _T_1462 ? 3'h4 : _GEN_4; // @[Conditional.scala 39:67:@22306.10]
  assign _GEN_6 = _T_1461 ? 3'h3 : _GEN_5; // @[Conditional.scala 39:67:@22301.8]
  assign _GEN_7 = _T_1460 ? 3'h2 : _GEN_6; // @[Conditional.scala 39:67:@22296.6]
  assign _GEN_8 = _T_1459 ? _GEN_0 : _GEN_7; // @[Conditional.scala 40:58:@22289.4]
  assign _T_1482 = state == 3'h0; // @[TensorAlu.scala 171:11:@22340.4]
  assign _T_1490 = _T_1441 & _T_1458; // @[TensorAlu.scala 173:31:@22347.4]
  assign _T_1491 = _T_1482 | _T_1490; // @[TensorAlu.scala 171:21:@22348.4]
  assign _T_1495 = uop_idx + 14'h1; // @[TensorAlu.scala 177:24:@22356.8]
  assign _T_1496 = uop_idx + 14'h1; // @[TensorAlu.scala 177:24:@22357.8]
  assign _GEN_9 = _T_1441 ? _T_1496 : uop_idx; // @[TensorAlu.scala 176:55:@22355.6]
  assign _T_1514 = _T_1490 & _T_1452; // @[TensorAlu.scala 187:33:@22378.6]
  assign _T_1516 = cnt_o + 14'h1; // @[TensorAlu.scala 189:20:@22380.8]
  assign _T_1517 = cnt_o + 14'h1; // @[TensorAlu.scala 189:20:@22381.8]
  assign _GEN_28 = {{3'd0}, dec_dst_0}; // @[TensorAlu.scala 190:20:@22383.8]
  assign _T_1518 = dst_o + _GEN_28; // @[TensorAlu.scala 190:20:@22383.8]
  assign _T_1519 = dst_o + _GEN_28; // @[TensorAlu.scala 190:20:@22384.8]
  assign _GEN_29 = {{3'd0}, dec_src_0}; // @[TensorAlu.scala 191:20:@22386.8]
  assign _T_1520 = src_o + _GEN_29; // @[TensorAlu.scala 191:20:@22386.8]
  assign _T_1521 = src_o + _GEN_29; // @[TensorAlu.scala 191:20:@22387.8]
  assign _GEN_11 = _T_1514 ? _T_1517 : cnt_o; // @[TensorAlu.scala 188:33:@22379.6]
  assign _GEN_12 = _T_1514 ? _T_1519 : dst_o; // @[TensorAlu.scala 188:33:@22379.6]
  assign _GEN_13 = _T_1514 ? _T_1521 : src_o; // @[TensorAlu.scala 188:33:@22379.6]
  assign _T_1526 = state == 3'h1; // @[TensorAlu.scala 198:20:@22397.6]
  assign _T_1527 = cnt_i == dec_lp_1; // @[TensorAlu.scala 198:42:@22398.6]
  assign _T_1528 = _T_1526 & _T_1527; // @[TensorAlu.scala 198:33:@22399.6]
  assign _T_1539 = cnt_i + 14'h1; // @[TensorAlu.scala 203:20:@22414.10]
  assign _T_1540 = cnt_i + 14'h1; // @[TensorAlu.scala 203:20:@22415.10]
  assign _GEN_30 = {{3'd0}, dec_dst_1}; // @[TensorAlu.scala 204:20:@22417.10]
  assign _T_1541 = dst_i + _GEN_30; // @[TensorAlu.scala 204:20:@22417.10]
  assign _T_1542 = dst_i + _GEN_30; // @[TensorAlu.scala 204:20:@22418.10]
  assign _GEN_31 = {{3'd0}, dec_src_1}; // @[TensorAlu.scala 205:20:@22420.10]
  assign _T_1543 = src_i + _GEN_31; // @[TensorAlu.scala 205:20:@22420.10]
  assign _T_1544 = src_i + _GEN_31; // @[TensorAlu.scala 205:20:@22421.10]
  assign _GEN_17 = _T_1490 ? _T_1540 : cnt_i; // @[TensorAlu.scala 202:84:@22413.8]
  assign _GEN_18 = _T_1490 ? _T_1542 : dst_i; // @[TensorAlu.scala 202:84:@22413.8]
  assign _GEN_19 = _T_1490 ? _T_1544 : src_i; // @[TensorAlu.scala 202:84:@22413.8]
  assign _GEN_20 = _T_1528 ? 14'h0 : _GEN_17; // @[TensorAlu.scala 198:56:@22400.6]
  assign _GEN_21 = _T_1528 ? dst_o : _GEN_18; // @[TensorAlu.scala 198:56:@22400.6]
  assign _GEN_22 = _T_1528 ? src_o : _GEN_19; // @[TensorAlu.scala 198:56:@22400.6]
  assign _T_1545 = state == 3'h2; // @[TensorAlu.scala 208:14:@22424.4]
  assign _T_1546 = _T_1545 & io_uop_data_valid; // @[TensorAlu.scala 208:30:@22425.4]
  assign _GEN_32 = {{3'd0}, io_uop_data_bits_u0}; // @[TensorAlu.scala 209:36:@22427.6]
  assign _T_1547 = _GEN_32 + dst_i; // @[TensorAlu.scala 209:36:@22427.6]
  assign _T_1548 = _GEN_32 + dst_i; // @[TensorAlu.scala 209:36:@22428.6]
  assign _GEN_33 = {{3'd0}, io_uop_data_bits_u1}; // @[TensorAlu.scala 210:36:@22430.6]
  assign _T_1549 = _GEN_33 + src_i; // @[TensorAlu.scala 210:36:@22430.6]
  assign _T_1550 = _GEN_33 + src_i; // @[TensorAlu.scala 210:36:@22431.6]
  assign _T_1552 = state == 3'h3; // @[TensorAlu.scala 218:32:@22437.4]
  assign _T_1553 = state == 3'h4; // @[TensorAlu.scala 218:58:@22438.4]
  assign _T_1554 = ~ dec_alu_use_imm; // @[TensorAlu.scala 218:77:@22439.4]
  assign _T_1555 = _T_1553 & _T_1554; // @[TensorAlu.scala 218:75:@22440.4]
  assign _T_1558 = _T_1552 ? uop_dst : uop_src; // @[TensorAlu.scala 219:28:@22444.4]
  assign _T_1863 = dec_alu_imm[15]; // @[TensorAlu.scala 226:27:@22449.4]
  assign _T_1866 = {16'hffff,dec_alu_imm}; // @[Cat.scala 30:58:@22451.4]
  assign tensorImm_data_bits_0_0 = _T_1863 ? _T_1866 : {{16'd0}, dec_alu_imm}; // @[TensorAlu.scala 226:15:@22452.4]
  assign _GEN_34 = {{1'd0}, dec_alu_op}; // @[TensorAlu.scala 232:26:@22529.4]
  assign isSHR = _GEN_34 == 3'h3; // @[TensorAlu.scala 232:26:@22529.4]
  assign neg_shift = isSHR & _T_1863; // @[TensorAlu.scala 233:25:@22531.4]
  assign _T_1945 = neg_shift ? 2'h0 : dec_alu_op; // @[TensorAlu.scala 234:40:@22532.4]
  assign _T_1949 = io_acc_rd_data_valid & _T_1440; // @[TensorAlu.scala 240:26:@22555.4]
  assign io_done = _T_1453 & _T_1458; // @[TensorAlu.scala 256:11:@22613.4]
  assign io_uop_idx_valid = state == 3'h1; // @[TensorAlu.scala 214:20:@22435.4]
  assign io_uop_idx_bits = uop_idx[10:0]; // @[TensorAlu.scala 215:19:@22436.4]
  assign io_acc_rd_idx_valid = _T_1552 | _T_1555; // @[TensorAlu.scala 218:23:@22442.4]
  assign io_acc_rd_idx_bits = _T_1558[10:0]; // @[TensorAlu.scala 219:22:@22445.4]
  assign io_acc_wr_valid = alu_io_acc_y_data_valid; // @[TensorAlu.scala 246:19:@22575.4]
  assign io_acc_wr_bits_idx = uop_dst[10:0]; // @[TensorAlu.scala 247:22:@22576.4]
  assign io_acc_wr_bits_data_0_0 = alu_io_acc_y_data_bits_0_0; // @[TensorAlu.scala 248:23:@22577.4]
  assign io_acc_wr_bits_data_0_1 = alu_io_acc_y_data_bits_0_1; // @[TensorAlu.scala 248:23:@22578.4]
  assign io_acc_wr_bits_data_0_2 = alu_io_acc_y_data_bits_0_2; // @[TensorAlu.scala 248:23:@22579.4]
  assign io_acc_wr_bits_data_0_3 = alu_io_acc_y_data_bits_0_3; // @[TensorAlu.scala 248:23:@22580.4]
  assign io_acc_wr_bits_data_0_4 = alu_io_acc_y_data_bits_0_4; // @[TensorAlu.scala 248:23:@22581.4]
  assign io_acc_wr_bits_data_0_5 = alu_io_acc_y_data_bits_0_5; // @[TensorAlu.scala 248:23:@22582.4]
  assign io_acc_wr_bits_data_0_6 = alu_io_acc_y_data_bits_0_6; // @[TensorAlu.scala 248:23:@22583.4]
  assign io_acc_wr_bits_data_0_7 = alu_io_acc_y_data_bits_0_7; // @[TensorAlu.scala 248:23:@22584.4]
  assign io_acc_wr_bits_data_0_8 = alu_io_acc_y_data_bits_0_8; // @[TensorAlu.scala 248:23:@22585.4]
  assign io_acc_wr_bits_data_0_9 = alu_io_acc_y_data_bits_0_9; // @[TensorAlu.scala 248:23:@22586.4]
  assign io_acc_wr_bits_data_0_10 = alu_io_acc_y_data_bits_0_10; // @[TensorAlu.scala 248:23:@22587.4]
  assign io_acc_wr_bits_data_0_11 = alu_io_acc_y_data_bits_0_11; // @[TensorAlu.scala 248:23:@22588.4]
  assign io_acc_wr_bits_data_0_12 = alu_io_acc_y_data_bits_0_12; // @[TensorAlu.scala 248:23:@22589.4]
  assign io_acc_wr_bits_data_0_13 = alu_io_acc_y_data_bits_0_13; // @[TensorAlu.scala 248:23:@22590.4]
  assign io_acc_wr_bits_data_0_14 = alu_io_acc_y_data_bits_0_14; // @[TensorAlu.scala 248:23:@22591.4]
  assign io_acc_wr_bits_data_0_15 = alu_io_acc_y_data_bits_0_15; // @[TensorAlu.scala 248:23:@22592.4]
  assign io_out_wr_valid = alu_io_out_data_valid; // @[TensorAlu.scala 251:19:@22593.4]
  assign io_out_wr_bits_idx = uop_dst[10:0]; // @[TensorAlu.scala 252:22:@22594.4]
  assign io_out_wr_bits_data_0_0 = alu_io_out_data_bits_0_0; // @[TensorAlu.scala 253:23:@22595.4]
  assign io_out_wr_bits_data_0_1 = alu_io_out_data_bits_0_1; // @[TensorAlu.scala 253:23:@22596.4]
  assign io_out_wr_bits_data_0_2 = alu_io_out_data_bits_0_2; // @[TensorAlu.scala 253:23:@22597.4]
  assign io_out_wr_bits_data_0_3 = alu_io_out_data_bits_0_3; // @[TensorAlu.scala 253:23:@22598.4]
  assign io_out_wr_bits_data_0_4 = alu_io_out_data_bits_0_4; // @[TensorAlu.scala 253:23:@22599.4]
  assign io_out_wr_bits_data_0_5 = alu_io_out_data_bits_0_5; // @[TensorAlu.scala 253:23:@22600.4]
  assign io_out_wr_bits_data_0_6 = alu_io_out_data_bits_0_6; // @[TensorAlu.scala 253:23:@22601.4]
  assign io_out_wr_bits_data_0_7 = alu_io_out_data_bits_0_7; // @[TensorAlu.scala 253:23:@22602.4]
  assign io_out_wr_bits_data_0_8 = alu_io_out_data_bits_0_8; // @[TensorAlu.scala 253:23:@22603.4]
  assign io_out_wr_bits_data_0_9 = alu_io_out_data_bits_0_9; // @[TensorAlu.scala 253:23:@22604.4]
  assign io_out_wr_bits_data_0_10 = alu_io_out_data_bits_0_10; // @[TensorAlu.scala 253:23:@22605.4]
  assign io_out_wr_bits_data_0_11 = alu_io_out_data_bits_0_11; // @[TensorAlu.scala 253:23:@22606.4]
  assign io_out_wr_bits_data_0_12 = alu_io_out_data_bits_0_12; // @[TensorAlu.scala 253:23:@22607.4]
  assign io_out_wr_bits_data_0_13 = alu_io_out_data_bits_0_13; // @[TensorAlu.scala 253:23:@22608.4]
  assign io_out_wr_bits_data_0_14 = alu_io_out_data_bits_0_14; // @[TensorAlu.scala 253:23:@22609.4]
  assign io_out_wr_bits_data_0_15 = alu_io_out_data_bits_0_15; // @[TensorAlu.scala 253:23:@22610.4]
  assign alu_clock = clock; // @[:@22219.4]
  assign alu_io_opcode = {neg_shift,_T_1945}; // @[TensorAlu.scala 235:17:@22534.4]
  assign alu_io_acc_a_data_valid = io_acc_rd_data_valid & _T_1553; // @[TensorAlu.scala 236:27:@22537.4]
  assign alu_io_acc_a_data_bits_0_0 = io_acc_rd_data_bits_0_0; // @[TensorAlu.scala 237:26:@22538.4]
  assign alu_io_acc_a_data_bits_0_1 = io_acc_rd_data_bits_0_1; // @[TensorAlu.scala 237:26:@22539.4]
  assign alu_io_acc_a_data_bits_0_2 = io_acc_rd_data_bits_0_2; // @[TensorAlu.scala 237:26:@22540.4]
  assign alu_io_acc_a_data_bits_0_3 = io_acc_rd_data_bits_0_3; // @[TensorAlu.scala 237:26:@22541.4]
  assign alu_io_acc_a_data_bits_0_4 = io_acc_rd_data_bits_0_4; // @[TensorAlu.scala 237:26:@22542.4]
  assign alu_io_acc_a_data_bits_0_5 = io_acc_rd_data_bits_0_5; // @[TensorAlu.scala 237:26:@22543.4]
  assign alu_io_acc_a_data_bits_0_6 = io_acc_rd_data_bits_0_6; // @[TensorAlu.scala 237:26:@22544.4]
  assign alu_io_acc_a_data_bits_0_7 = io_acc_rd_data_bits_0_7; // @[TensorAlu.scala 237:26:@22545.4]
  assign alu_io_acc_a_data_bits_0_8 = io_acc_rd_data_bits_0_8; // @[TensorAlu.scala 237:26:@22546.4]
  assign alu_io_acc_a_data_bits_0_9 = io_acc_rd_data_bits_0_9; // @[TensorAlu.scala 237:26:@22547.4]
  assign alu_io_acc_a_data_bits_0_10 = io_acc_rd_data_bits_0_10; // @[TensorAlu.scala 237:26:@22548.4]
  assign alu_io_acc_a_data_bits_0_11 = io_acc_rd_data_bits_0_11; // @[TensorAlu.scala 237:26:@22549.4]
  assign alu_io_acc_a_data_bits_0_12 = io_acc_rd_data_bits_0_12; // @[TensorAlu.scala 237:26:@22550.4]
  assign alu_io_acc_a_data_bits_0_13 = io_acc_rd_data_bits_0_13; // @[TensorAlu.scala 237:26:@22551.4]
  assign alu_io_acc_a_data_bits_0_14 = io_acc_rd_data_bits_0_14; // @[TensorAlu.scala 237:26:@22552.4]
  assign alu_io_acc_a_data_bits_0_15 = io_acc_rd_data_bits_0_15; // @[TensorAlu.scala 237:26:@22553.4]
  assign alu_io_acc_b_data_valid = dec_alu_use_imm ? _T_1553 : _T_1949; // @[TensorAlu.scala 238:27:@22557.4]
  assign alu_io_acc_b_data_bits_0_0 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_0; // @[TensorAlu.scala 241:26:@22559.4]
  assign alu_io_acc_b_data_bits_0_1 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_1; // @[TensorAlu.scala 241:26:@22560.4]
  assign alu_io_acc_b_data_bits_0_2 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_2; // @[TensorAlu.scala 241:26:@22561.4]
  assign alu_io_acc_b_data_bits_0_3 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_3; // @[TensorAlu.scala 241:26:@22562.4]
  assign alu_io_acc_b_data_bits_0_4 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_4; // @[TensorAlu.scala 241:26:@22563.4]
  assign alu_io_acc_b_data_bits_0_5 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_5; // @[TensorAlu.scala 241:26:@22564.4]
  assign alu_io_acc_b_data_bits_0_6 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_6; // @[TensorAlu.scala 241:26:@22565.4]
  assign alu_io_acc_b_data_bits_0_7 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_7; // @[TensorAlu.scala 241:26:@22566.4]
  assign alu_io_acc_b_data_bits_0_8 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_8; // @[TensorAlu.scala 241:26:@22567.4]
  assign alu_io_acc_b_data_bits_0_9 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_9; // @[TensorAlu.scala 241:26:@22568.4]
  assign alu_io_acc_b_data_bits_0_10 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_10; // @[TensorAlu.scala 241:26:@22569.4]
  assign alu_io_acc_b_data_bits_0_11 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_11; // @[TensorAlu.scala 241:26:@22570.4]
  assign alu_io_acc_b_data_bits_0_12 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_12; // @[TensorAlu.scala 241:26:@22571.4]
  assign alu_io_acc_b_data_bits_0_13 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_13; // @[TensorAlu.scala 241:26:@22572.4]
  assign alu_io_acc_b_data_bits_0_14 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_14; // @[TensorAlu.scala 241:26:@22573.4]
  assign alu_io_acc_b_data_bits_0_15 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_15; // @[TensorAlu.scala 241:26:@22574.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  uop_idx = _RAND_1[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  uop_dst = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  uop_src = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cnt_o = _RAND_4[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  dst_o = _RAND_5[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  src_o = _RAND_6[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  cnt_i = _RAND_7[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  dst_i = _RAND_8[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  src_i = _RAND_9[13:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_1459) begin
        if (io_start) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_1460) begin
          state <= 3'h2;
        end else begin
          if (_T_1461) begin
            state <= 3'h3;
          end else begin
            if (_T_1462) begin
              state <= 3'h4;
            end else begin
              if (_T_1463) begin
                state <= 3'h5;
              end else begin
                if (_T_1464) begin
                  if (alu_io_out_data_valid) begin
                    if (_T_1481) begin
                      state <= 3'h0;
                    end else begin
                      state <= 3'h1;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_1491) begin
      uop_idx <= {{1'd0}, dec_uop_begin};
    end else begin
      if (_T_1441) begin
        uop_idx <= _T_1496;
      end
    end
    if (_T_1546) begin
      uop_dst <= _T_1548;
    end
    if (_T_1546) begin
      uop_src <= _T_1550;
    end
    if (_T_1482) begin
      cnt_o <= 14'h0;
    end else begin
      if (_T_1514) begin
        cnt_o <= _T_1517;
      end
    end
    if (_T_1482) begin
      dst_o <= 14'h0;
    end else begin
      if (_T_1514) begin
        dst_o <= _T_1519;
      end
    end
    if (_T_1482) begin
      src_o <= 14'h0;
    end else begin
      if (_T_1514) begin
        src_o <= _T_1521;
      end
    end
    if (_T_1482) begin
      cnt_i <= 14'h0;
    end else begin
      if (_T_1528) begin
        cnt_i <= 14'h0;
      end else begin
        if (_T_1490) begin
          cnt_i <= _T_1540;
        end
      end
    end
    if (_T_1482) begin
      dst_i <= 14'h0;
    end else begin
      if (_T_1528) begin
        dst_i <= dst_o;
      end else begin
        if (_T_1490) begin
          dst_i <= _T_1542;
        end
      end
    end
    if (_T_1482) begin
      src_i <= 14'h0;
    end else begin
      if (_T_1528) begin
        src_i <= src_o;
      end else begin
        if (_T_1490) begin
          src_i <= _T_1544;
        end
      end
    end
  end
endmodule
module ComputeDecode( // @[:@22666.2]
  input  [127:0] io_inst, // @[:@22669.4]
  output         io_push_next, // @[:@22669.4]
  output         io_push_prev, // @[:@22669.4]
  output         io_pop_next, // @[:@22669.4]
  output         io_pop_prev, // @[:@22669.4]
  output         io_isLoadAcc, // @[:@22669.4]
  output         io_isLoadUop, // @[:@22669.4]
  output         io_isSync, // @[:@22669.4]
  output         io_isAlu, // @[:@22669.4]
  output         io_isGemm, // @[:@22669.4]
  output         io_isFinish // @[:@22669.4]
);
  wire [15:0] dec_xsize; // @[Decode.scala 200:29:@22694.4]
  wire [127:0] _T_49; // @[Decode.scala 205:27:@22710.4]
  wire  _T_50; // @[Decode.scala 205:27:@22711.4]
  wire  _T_52; // @[Decode.scala 205:48:@22712.4]
  wire  _T_57; // @[Decode.scala 206:27:@22716.4]
  wire  _T_69; // @[Decode.scala 207:34:@22724.4]
  wire  _T_71; // @[Decode.scala 207:66:@22725.4]
  wire [127:0] _T_75; // @[Decode.scala 208:23:@22728.4]
  wire  _T_76; // @[Decode.scala 208:23:@22729.4]
  wire  _T_80; // @[Decode.scala 208:42:@22731.4]
  wire  _T_81; // @[Decode.scala 208:32:@22732.4]
  wire  _T_85; // @[Decode.scala 208:61:@22734.4]
  wire  _T_86; // @[Decode.scala 208:51:@22735.4]
  wire  _T_90; // @[Decode.scala 208:80:@22737.4]
  wire [127:0] _T_94; // @[Decode.scala 209:24:@22740.4]
  assign dec_xsize = io_inst[95:80]; // @[Decode.scala 200:29:@22694.4]
  assign _T_49 = io_inst & 128'h187; // @[Decode.scala 205:27:@22710.4]
  assign _T_50 = 128'h180 == _T_49; // @[Decode.scala 205:27:@22711.4]
  assign _T_52 = dec_xsize != 16'h0; // @[Decode.scala 205:48:@22712.4]
  assign _T_57 = 128'h0 == _T_49; // @[Decode.scala 206:27:@22716.4]
  assign _T_69 = _T_50 | _T_57; // @[Decode.scala 207:34:@22724.4]
  assign _T_71 = dec_xsize == 16'h0; // @[Decode.scala 207:66:@22725.4]
  assign _T_75 = io_inst & 128'h3000000000000000000000000007; // @[Decode.scala 208:23:@22728.4]
  assign _T_76 = 128'h4 == _T_75; // @[Decode.scala 208:23:@22729.4]
  assign _T_80 = 128'h1000000000000000000000000004 == _T_75; // @[Decode.scala 208:42:@22731.4]
  assign _T_81 = _T_76 | _T_80; // @[Decode.scala 208:32:@22732.4]
  assign _T_85 = 128'h2000000000000000000000000004 == _T_75; // @[Decode.scala 208:61:@22734.4]
  assign _T_86 = _T_81 | _T_85; // @[Decode.scala 208:51:@22735.4]
  assign _T_90 = 128'h3000000000000000000000000004 == _T_75; // @[Decode.scala 208:80:@22737.4]
  assign _T_94 = io_inst & 128'h7; // @[Decode.scala 209:24:@22740.4]
  assign io_push_next = io_inst[6]; // @[Decode.scala 201:16:@22706.4]
  assign io_push_prev = io_inst[5]; // @[Decode.scala 202:16:@22707.4]
  assign io_pop_next = io_inst[4]; // @[Decode.scala 203:15:@22708.4]
  assign io_pop_prev = io_inst[3]; // @[Decode.scala 204:15:@22709.4]
  assign io_isLoadAcc = _T_50 & _T_52; // @[Decode.scala 205:16:@22714.4]
  assign io_isLoadUop = _T_57 & _T_52; // @[Decode.scala 206:16:@22719.4]
  assign io_isSync = _T_69 & _T_71; // @[Decode.scala 207:13:@22727.4]
  assign io_isAlu = _T_86 | _T_90; // @[Decode.scala 208:12:@22739.4]
  assign io_isGemm = 128'h2 == _T_94; // @[Decode.scala 209:13:@22742.4]
  assign io_isFinish = 128'h3 == _T_94; // @[Decode.scala 210:15:@22745.4]
endmodule
module Compute( // @[:@22747.2]
  input          clock, // @[:@22748.4]
  input          reset, // @[:@22749.4]
  input          io_i_post_0, // @[:@22750.4]
  input          io_i_post_1, // @[:@22750.4]
  output         io_o_post_0, // @[:@22750.4]
  output         io_o_post_1, // @[:@22750.4]
  output         io_inst_ready, // @[:@22750.4]
  input          io_inst_valid, // @[:@22750.4]
  input  [127:0] io_inst_bits, // @[:@22750.4]
  input  [31:0]  io_uop_baddr, // @[:@22750.4]
  input  [31:0]  io_acc_baddr, // @[:@22750.4]
  input          io_vme_rd_0_cmd_ready, // @[:@22750.4]
  output         io_vme_rd_0_cmd_valid, // @[:@22750.4]
  output [31:0]  io_vme_rd_0_cmd_bits_addr, // @[:@22750.4]
  output [7:0]   io_vme_rd_0_cmd_bits_len, // @[:@22750.4]
  output         io_vme_rd_0_data_ready, // @[:@22750.4]
  input          io_vme_rd_0_data_valid, // @[:@22750.4]
  input  [63:0]  io_vme_rd_0_data_bits, // @[:@22750.4]
  input          io_vme_rd_1_cmd_ready, // @[:@22750.4]
  output         io_vme_rd_1_cmd_valid, // @[:@22750.4]
  output [31:0]  io_vme_rd_1_cmd_bits_addr, // @[:@22750.4]
  output [7:0]   io_vme_rd_1_cmd_bits_len, // @[:@22750.4]
  output         io_vme_rd_1_data_ready, // @[:@22750.4]
  input          io_vme_rd_1_data_valid, // @[:@22750.4]
  input  [63:0]  io_vme_rd_1_data_bits, // @[:@22750.4]
  output         io_inp_rd_idx_valid, // @[:@22750.4]
  output [10:0]  io_inp_rd_idx_bits, // @[:@22750.4]
  input          io_inp_rd_data_valid, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_0, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_1, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_2, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_3, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_4, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_5, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_6, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_7, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_8, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_9, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_10, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_11, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_12, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_13, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_14, // @[:@22750.4]
  input  [7:0]   io_inp_rd_data_bits_0_15, // @[:@22750.4]
  output         io_wgt_rd_idx_valid, // @[:@22750.4]
  output [9:0]   io_wgt_rd_idx_bits, // @[:@22750.4]
  input          io_wgt_rd_data_valid, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_0_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_1_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_2_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_3_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_4_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_5_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_6_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_7_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_8_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_9_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_10_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_11_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_12_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_13_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_14_15, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_0, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_1, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_2, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_3, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_4, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_5, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_6, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_7, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_8, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_9, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_10, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_11, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_12, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_13, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_14, // @[:@22750.4]
  input  [7:0]   io_wgt_rd_data_bits_15_15, // @[:@22750.4]
  output         io_out_wr_valid, // @[:@22750.4]
  output [10:0]  io_out_wr_bits_idx, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_0, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_1, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_2, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_3, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_4, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_5, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_6, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_7, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_8, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_9, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_10, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_11, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_12, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_13, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_14, // @[:@22750.4]
  output [7:0]   io_out_wr_bits_data_0_15, // @[:@22750.4]
  output         io_finish, // @[:@22750.4]
  output         io_acc_wr_event // @[:@22750.4]
);
  wire  s_0_clock; // @[Compute.scala 54:11:@22753.4]
  wire  s_0_reset; // @[Compute.scala 54:11:@22753.4]
  wire  s_0_io_spost; // @[Compute.scala 54:11:@22753.4]
  wire  s_0_io_swait; // @[Compute.scala 54:11:@22753.4]
  wire  s_0_io_sready; // @[Compute.scala 54:11:@22753.4]
  wire  s_1_clock; // @[Compute.scala 54:11:@22756.4]
  wire  s_1_reset; // @[Compute.scala 54:11:@22756.4]
  wire  s_1_io_spost; // @[Compute.scala 54:11:@22756.4]
  wire  s_1_io_swait; // @[Compute.scala 54:11:@22756.4]
  wire  s_1_io_sready; // @[Compute.scala 54:11:@22756.4]
  wire  loadUop_clock; // @[Compute.scala 56:23:@22759.4]
  wire  loadUop_reset; // @[Compute.scala 56:23:@22759.4]
  wire  loadUop_io_start; // @[Compute.scala 56:23:@22759.4]
  wire  loadUop_io_done; // @[Compute.scala 56:23:@22759.4]
  wire [127:0] loadUop_io_inst; // @[Compute.scala 56:23:@22759.4]
  wire [31:0] loadUop_io_baddr; // @[Compute.scala 56:23:@22759.4]
  wire  loadUop_io_vme_rd_cmd_ready; // @[Compute.scala 56:23:@22759.4]
  wire  loadUop_io_vme_rd_cmd_valid; // @[Compute.scala 56:23:@22759.4]
  wire [31:0] loadUop_io_vme_rd_cmd_bits_addr; // @[Compute.scala 56:23:@22759.4]
  wire [7:0] loadUop_io_vme_rd_cmd_bits_len; // @[Compute.scala 56:23:@22759.4]
  wire  loadUop_io_vme_rd_data_ready; // @[Compute.scala 56:23:@22759.4]
  wire  loadUop_io_vme_rd_data_valid; // @[Compute.scala 56:23:@22759.4]
  wire [63:0] loadUop_io_vme_rd_data_bits; // @[Compute.scala 56:23:@22759.4]
  wire  loadUop_io_uop_idx_valid; // @[Compute.scala 56:23:@22759.4]
  wire [10:0] loadUop_io_uop_idx_bits; // @[Compute.scala 56:23:@22759.4]
  wire  loadUop_io_uop_data_valid; // @[Compute.scala 56:23:@22759.4]
  wire [9:0] loadUop_io_uop_data_bits_u2; // @[Compute.scala 56:23:@22759.4]
  wire [10:0] loadUop_io_uop_data_bits_u1; // @[Compute.scala 56:23:@22759.4]
  wire [10:0] loadUop_io_uop_data_bits_u0; // @[Compute.scala 56:23:@22759.4]
  wire  tensorAcc_clock; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_reset; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_io_start; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_io_done; // @[Compute.scala 57:25:@22762.4]
  wire [127:0] tensorAcc_io_inst; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_baddr; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_io_vme_rd_cmd_ready; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_io_vme_rd_cmd_valid; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_vme_rd_cmd_bits_addr; // @[Compute.scala 57:25:@22762.4]
  wire [7:0] tensorAcc_io_vme_rd_cmd_bits_len; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_io_vme_rd_data_ready; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_io_vme_rd_data_valid; // @[Compute.scala 57:25:@22762.4]
  wire [63:0] tensorAcc_io_vme_rd_data_bits; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_io_tensor_rd_idx_valid; // @[Compute.scala 57:25:@22762.4]
  wire [10:0] tensorAcc_io_tensor_rd_idx_bits; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_io_tensor_rd_data_valid; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_0; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_1; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_2; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_3; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_4; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_5; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_6; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_7; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_8; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_9; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_10; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_11; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_12; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_13; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_14; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_15; // @[Compute.scala 57:25:@22762.4]
  wire  tensorAcc_io_tensor_wr_valid; // @[Compute.scala 57:25:@22762.4]
  wire [10:0] tensorAcc_io_tensor_wr_bits_idx; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_0; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_1; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_2; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_3; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_4; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_5; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_6; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_7; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_8; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_9; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_10; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_11; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_12; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_13; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_14; // @[Compute.scala 57:25:@22762.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_15; // @[Compute.scala 57:25:@22762.4]
  wire  tensorGemm_clock; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_reset; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_start; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_done; // @[Compute.scala 58:26:@22765.4]
  wire [127:0] tensorGemm_io_inst; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_uop_idx_valid; // @[Compute.scala 58:26:@22765.4]
  wire [10:0] tensorGemm_io_uop_idx_bits; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_uop_data_valid; // @[Compute.scala 58:26:@22765.4]
  wire [9:0] tensorGemm_io_uop_data_bits_u2; // @[Compute.scala 58:26:@22765.4]
  wire [10:0] tensorGemm_io_uop_data_bits_u1; // @[Compute.scala 58:26:@22765.4]
  wire [10:0] tensorGemm_io_uop_data_bits_u0; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_inp_rd_idx_valid; // @[Compute.scala 58:26:@22765.4]
  wire [10:0] tensorGemm_io_inp_rd_idx_bits; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_inp_rd_data_valid; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_15; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_wgt_rd_idx_valid; // @[Compute.scala 58:26:@22765.4]
  wire [9:0] tensorGemm_io_wgt_rd_idx_bits; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_wgt_rd_data_valid; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_15; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_15; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_acc_rd_idx_valid; // @[Compute.scala 58:26:@22765.4]
  wire [10:0] tensorGemm_io_acc_rd_idx_bits; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_acc_rd_data_valid; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_0; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_1; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_2; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_3; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_4; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_5; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_6; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_7; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_8; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_9; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_10; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_11; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_12; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_13; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_14; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_15; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_acc_wr_valid; // @[Compute.scala 58:26:@22765.4]
  wire [10:0] tensorGemm_io_acc_wr_bits_idx; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_0; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_1; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_2; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_3; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_4; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_5; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_6; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_7; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_8; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_9; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_10; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_11; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_12; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_13; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_14; // @[Compute.scala 58:26:@22765.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_15; // @[Compute.scala 58:26:@22765.4]
  wire  tensorGemm_io_out_wr_valid; // @[Compute.scala 58:26:@22765.4]
  wire [10:0] tensorGemm_io_out_wr_bits_idx; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_0; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_1; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_2; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_3; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_4; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_5; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_6; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_7; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_8; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_9; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_10; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_11; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_12; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_13; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_14; // @[Compute.scala 58:26:@22765.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_15; // @[Compute.scala 58:26:@22765.4]
  wire  tensorAlu_clock; // @[Compute.scala 59:25:@22768.4]
  wire  tensorAlu_reset; // @[Compute.scala 59:25:@22768.4]
  wire  tensorAlu_io_start; // @[Compute.scala 59:25:@22768.4]
  wire  tensorAlu_io_done; // @[Compute.scala 59:25:@22768.4]
  wire [127:0] tensorAlu_io_inst; // @[Compute.scala 59:25:@22768.4]
  wire  tensorAlu_io_uop_idx_valid; // @[Compute.scala 59:25:@22768.4]
  wire [10:0] tensorAlu_io_uop_idx_bits; // @[Compute.scala 59:25:@22768.4]
  wire  tensorAlu_io_uop_data_valid; // @[Compute.scala 59:25:@22768.4]
  wire [10:0] tensorAlu_io_uop_data_bits_u1; // @[Compute.scala 59:25:@22768.4]
  wire [10:0] tensorAlu_io_uop_data_bits_u0; // @[Compute.scala 59:25:@22768.4]
  wire  tensorAlu_io_acc_rd_idx_valid; // @[Compute.scala 59:25:@22768.4]
  wire [10:0] tensorAlu_io_acc_rd_idx_bits; // @[Compute.scala 59:25:@22768.4]
  wire  tensorAlu_io_acc_rd_data_valid; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_0; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_1; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_2; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_3; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_4; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_5; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_6; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_7; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_8; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_9; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_10; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_11; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_12; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_13; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_14; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_15; // @[Compute.scala 59:25:@22768.4]
  wire  tensorAlu_io_acc_wr_valid; // @[Compute.scala 59:25:@22768.4]
  wire [10:0] tensorAlu_io_acc_wr_bits_idx; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_0; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_1; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_2; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_3; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_4; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_5; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_6; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_7; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_8; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_9; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_10; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_11; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_12; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_13; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_14; // @[Compute.scala 59:25:@22768.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_15; // @[Compute.scala 59:25:@22768.4]
  wire  tensorAlu_io_out_wr_valid; // @[Compute.scala 59:25:@22768.4]
  wire [10:0] tensorAlu_io_out_wr_bits_idx; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_0; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_1; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_2; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_3; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_4; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_5; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_6; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_7; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_8; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_9; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_10; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_11; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_12; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_13; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_14; // @[Compute.scala 59:25:@22768.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_15; // @[Compute.scala 59:25:@22768.4]
  wire  inst_q_clock; // @[Compute.scala 61:22:@22771.4]
  wire  inst_q_reset; // @[Compute.scala 61:22:@22771.4]
  wire  inst_q_io_enq_ready; // @[Compute.scala 61:22:@22771.4]
  wire  inst_q_io_enq_valid; // @[Compute.scala 61:22:@22771.4]
  wire [127:0] inst_q_io_enq_bits; // @[Compute.scala 61:22:@22771.4]
  wire  inst_q_io_deq_ready; // @[Compute.scala 61:22:@22771.4]
  wire  inst_q_io_deq_valid; // @[Compute.scala 61:22:@22771.4]
  wire [127:0] inst_q_io_deq_bits; // @[Compute.scala 61:22:@22771.4]
  wire [127:0] dec_io_inst; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_push_next; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_push_prev; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_pop_next; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_pop_prev; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_isLoadAcc; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_isLoadUop; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_isSync; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_isAlu; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_isGemm; // @[Compute.scala 64:19:@22774.4]
  wire  dec_io_isFinish; // @[Compute.scala 64:19:@22774.4]
  reg [1:0] state; // @[Compute.scala 51:22:@22752.4]
  reg [31:0] _RAND_0;
  wire [4:0] inst_type; // @[Cat.scala 30:58:@22781.4]
  wire  _T_7054; // @[Compute.scala 74:40:@22782.4]
  wire  sprev; // @[Compute.scala 74:35:@22783.4]
  wire  _T_7056; // @[Compute.scala 75:40:@22784.4]
  wire  snext; // @[Compute.scala 75:35:@22785.4]
  wire  start; // @[Compute.scala 76:21:@22786.4]
  wire  _T_7064; // @[Mux.scala 46:19:@22787.4]
  wire  _T_7066; // @[Mux.scala 46:19:@22789.4]
  wire  _T_7067; // @[Mux.scala 46:16:@22790.4]
  wire  _T_7068; // @[Mux.scala 46:19:@22791.4]
  wire  _T_7069; // @[Mux.scala 46:16:@22792.4]
  wire  _T_7070; // @[Mux.scala 46:19:@22793.4]
  wire  _T_7071; // @[Mux.scala 46:16:@22794.4]
  wire  _T_7072; // @[Mux.scala 46:19:@22795.4]
  wire  done; // @[Mux.scala 46:16:@22796.4]
  wire  _T_7073; // @[Conditional.scala 37:30:@22797.4]
  wire  _T_7075; // @[Compute.scala 96:30:@22804.10]
  wire [1:0] _GEN_0; // @[Compute.scala 96:35:@22805.10]
  wire [1:0] _GEN_1; // @[Compute.scala 94:29:@22800.8]
  wire [1:0] _GEN_2; // @[Compute.scala 93:19:@22799.6]
  wire  _T_7076; // @[Conditional.scala 37:30:@22811.6]
  wire  _T_7077; // @[Conditional.scala 37:30:@22816.8]
  wire [1:0] _GEN_3; // @[Compute.scala 105:18:@22818.10]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@22817.8]
  wire [1:0] _GEN_5; // @[Conditional.scala 39:67:@22812.6]
  wire [1:0] _GEN_6; // @[Conditional.scala 40:58:@22798.4]
  wire  _T_7078; // @[Compute.scala 113:33:@22825.4]
  wire  _T_7079; // @[Compute.scala 113:42:@22826.4]
  wire  _T_7080; // @[Compute.scala 113:59:@22827.4]
  wire  _T_7081; // @[Compute.scala 113:50:@22828.4]
  wire  _T_7082; // @[Compute.scala 116:29:@22830.4]
  wire  _T_7083; // @[Compute.scala 116:39:@22831.4]
  Semaphore s_0 ( // @[Compute.scala 54:11:@22753.4]
    .clock(s_0_clock),
    .reset(s_0_reset),
    .io_spost(s_0_io_spost),
    .io_swait(s_0_io_swait),
    .io_sready(s_0_io_sready)
  );
  Semaphore s_1 ( // @[Compute.scala 54:11:@22756.4]
    .clock(s_1_clock),
    .reset(s_1_reset),
    .io_spost(s_1_io_spost),
    .io_swait(s_1_io_swait),
    .io_sready(s_1_io_sready)
  );
  LoadUop loadUop ( // @[Compute.scala 56:23:@22759.4]
    .clock(loadUop_clock),
    .reset(loadUop_reset),
    .io_start(loadUop_io_start),
    .io_done(loadUop_io_done),
    .io_inst(loadUop_io_inst),
    .io_baddr(loadUop_io_baddr),
    .io_vme_rd_cmd_ready(loadUop_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(loadUop_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(loadUop_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(loadUop_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(loadUop_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(loadUop_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(loadUop_io_vme_rd_data_bits),
    .io_uop_idx_valid(loadUop_io_uop_idx_valid),
    .io_uop_idx_bits(loadUop_io_uop_idx_bits),
    .io_uop_data_valid(loadUop_io_uop_data_valid),
    .io_uop_data_bits_u2(loadUop_io_uop_data_bits_u2),
    .io_uop_data_bits_u1(loadUop_io_uop_data_bits_u1),
    .io_uop_data_bits_u0(loadUop_io_uop_data_bits_u0)
  );
  TensorLoad_2 tensorAcc ( // @[Compute.scala 57:25:@22762.4]
    .clock(tensorAcc_clock),
    .reset(tensorAcc_reset),
    .io_start(tensorAcc_io_start),
    .io_done(tensorAcc_io_done),
    .io_inst(tensorAcc_io_inst),
    .io_baddr(tensorAcc_io_baddr),
    .io_vme_rd_cmd_ready(tensorAcc_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorAcc_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorAcc_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorAcc_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(tensorAcc_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorAcc_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(tensorAcc_io_vme_rd_data_bits),
    .io_tensor_rd_idx_valid(tensorAcc_io_tensor_rd_idx_valid),
    .io_tensor_rd_idx_bits(tensorAcc_io_tensor_rd_idx_bits),
    .io_tensor_rd_data_valid(tensorAcc_io_tensor_rd_data_valid),
    .io_tensor_rd_data_bits_0_0(tensorAcc_io_tensor_rd_data_bits_0_0),
    .io_tensor_rd_data_bits_0_1(tensorAcc_io_tensor_rd_data_bits_0_1),
    .io_tensor_rd_data_bits_0_2(tensorAcc_io_tensor_rd_data_bits_0_2),
    .io_tensor_rd_data_bits_0_3(tensorAcc_io_tensor_rd_data_bits_0_3),
    .io_tensor_rd_data_bits_0_4(tensorAcc_io_tensor_rd_data_bits_0_4),
    .io_tensor_rd_data_bits_0_5(tensorAcc_io_tensor_rd_data_bits_0_5),
    .io_tensor_rd_data_bits_0_6(tensorAcc_io_tensor_rd_data_bits_0_6),
    .io_tensor_rd_data_bits_0_7(tensorAcc_io_tensor_rd_data_bits_0_7),
    .io_tensor_rd_data_bits_0_8(tensorAcc_io_tensor_rd_data_bits_0_8),
    .io_tensor_rd_data_bits_0_9(tensorAcc_io_tensor_rd_data_bits_0_9),
    .io_tensor_rd_data_bits_0_10(tensorAcc_io_tensor_rd_data_bits_0_10),
    .io_tensor_rd_data_bits_0_11(tensorAcc_io_tensor_rd_data_bits_0_11),
    .io_tensor_rd_data_bits_0_12(tensorAcc_io_tensor_rd_data_bits_0_12),
    .io_tensor_rd_data_bits_0_13(tensorAcc_io_tensor_rd_data_bits_0_13),
    .io_tensor_rd_data_bits_0_14(tensorAcc_io_tensor_rd_data_bits_0_14),
    .io_tensor_rd_data_bits_0_15(tensorAcc_io_tensor_rd_data_bits_0_15),
    .io_tensor_wr_valid(tensorAcc_io_tensor_wr_valid),
    .io_tensor_wr_bits_idx(tensorAcc_io_tensor_wr_bits_idx),
    .io_tensor_wr_bits_data_0_0(tensorAcc_io_tensor_wr_bits_data_0_0),
    .io_tensor_wr_bits_data_0_1(tensorAcc_io_tensor_wr_bits_data_0_1),
    .io_tensor_wr_bits_data_0_2(tensorAcc_io_tensor_wr_bits_data_0_2),
    .io_tensor_wr_bits_data_0_3(tensorAcc_io_tensor_wr_bits_data_0_3),
    .io_tensor_wr_bits_data_0_4(tensorAcc_io_tensor_wr_bits_data_0_4),
    .io_tensor_wr_bits_data_0_5(tensorAcc_io_tensor_wr_bits_data_0_5),
    .io_tensor_wr_bits_data_0_6(tensorAcc_io_tensor_wr_bits_data_0_6),
    .io_tensor_wr_bits_data_0_7(tensorAcc_io_tensor_wr_bits_data_0_7),
    .io_tensor_wr_bits_data_0_8(tensorAcc_io_tensor_wr_bits_data_0_8),
    .io_tensor_wr_bits_data_0_9(tensorAcc_io_tensor_wr_bits_data_0_9),
    .io_tensor_wr_bits_data_0_10(tensorAcc_io_tensor_wr_bits_data_0_10),
    .io_tensor_wr_bits_data_0_11(tensorAcc_io_tensor_wr_bits_data_0_11),
    .io_tensor_wr_bits_data_0_12(tensorAcc_io_tensor_wr_bits_data_0_12),
    .io_tensor_wr_bits_data_0_13(tensorAcc_io_tensor_wr_bits_data_0_13),
    .io_tensor_wr_bits_data_0_14(tensorAcc_io_tensor_wr_bits_data_0_14),
    .io_tensor_wr_bits_data_0_15(tensorAcc_io_tensor_wr_bits_data_0_15)
  );
  TensorGemm tensorGemm ( // @[Compute.scala 58:26:@22765.4]
    .clock(tensorGemm_clock),
    .reset(tensorGemm_reset),
    .io_start(tensorGemm_io_start),
    .io_done(tensorGemm_io_done),
    .io_inst(tensorGemm_io_inst),
    .io_uop_idx_valid(tensorGemm_io_uop_idx_valid),
    .io_uop_idx_bits(tensorGemm_io_uop_idx_bits),
    .io_uop_data_valid(tensorGemm_io_uop_data_valid),
    .io_uop_data_bits_u2(tensorGemm_io_uop_data_bits_u2),
    .io_uop_data_bits_u1(tensorGemm_io_uop_data_bits_u1),
    .io_uop_data_bits_u0(tensorGemm_io_uop_data_bits_u0),
    .io_inp_rd_idx_valid(tensorGemm_io_inp_rd_idx_valid),
    .io_inp_rd_idx_bits(tensorGemm_io_inp_rd_idx_bits),
    .io_inp_rd_data_valid(tensorGemm_io_inp_rd_data_valid),
    .io_inp_rd_data_bits_0_0(tensorGemm_io_inp_rd_data_bits_0_0),
    .io_inp_rd_data_bits_0_1(tensorGemm_io_inp_rd_data_bits_0_1),
    .io_inp_rd_data_bits_0_2(tensorGemm_io_inp_rd_data_bits_0_2),
    .io_inp_rd_data_bits_0_3(tensorGemm_io_inp_rd_data_bits_0_3),
    .io_inp_rd_data_bits_0_4(tensorGemm_io_inp_rd_data_bits_0_4),
    .io_inp_rd_data_bits_0_5(tensorGemm_io_inp_rd_data_bits_0_5),
    .io_inp_rd_data_bits_0_6(tensorGemm_io_inp_rd_data_bits_0_6),
    .io_inp_rd_data_bits_0_7(tensorGemm_io_inp_rd_data_bits_0_7),
    .io_inp_rd_data_bits_0_8(tensorGemm_io_inp_rd_data_bits_0_8),
    .io_inp_rd_data_bits_0_9(tensorGemm_io_inp_rd_data_bits_0_9),
    .io_inp_rd_data_bits_0_10(tensorGemm_io_inp_rd_data_bits_0_10),
    .io_inp_rd_data_bits_0_11(tensorGemm_io_inp_rd_data_bits_0_11),
    .io_inp_rd_data_bits_0_12(tensorGemm_io_inp_rd_data_bits_0_12),
    .io_inp_rd_data_bits_0_13(tensorGemm_io_inp_rd_data_bits_0_13),
    .io_inp_rd_data_bits_0_14(tensorGemm_io_inp_rd_data_bits_0_14),
    .io_inp_rd_data_bits_0_15(tensorGemm_io_inp_rd_data_bits_0_15),
    .io_wgt_rd_idx_valid(tensorGemm_io_wgt_rd_idx_valid),
    .io_wgt_rd_idx_bits(tensorGemm_io_wgt_rd_idx_bits),
    .io_wgt_rd_data_valid(tensorGemm_io_wgt_rd_data_valid),
    .io_wgt_rd_data_bits_0_0(tensorGemm_io_wgt_rd_data_bits_0_0),
    .io_wgt_rd_data_bits_0_1(tensorGemm_io_wgt_rd_data_bits_0_1),
    .io_wgt_rd_data_bits_0_2(tensorGemm_io_wgt_rd_data_bits_0_2),
    .io_wgt_rd_data_bits_0_3(tensorGemm_io_wgt_rd_data_bits_0_3),
    .io_wgt_rd_data_bits_0_4(tensorGemm_io_wgt_rd_data_bits_0_4),
    .io_wgt_rd_data_bits_0_5(tensorGemm_io_wgt_rd_data_bits_0_5),
    .io_wgt_rd_data_bits_0_6(tensorGemm_io_wgt_rd_data_bits_0_6),
    .io_wgt_rd_data_bits_0_7(tensorGemm_io_wgt_rd_data_bits_0_7),
    .io_wgt_rd_data_bits_0_8(tensorGemm_io_wgt_rd_data_bits_0_8),
    .io_wgt_rd_data_bits_0_9(tensorGemm_io_wgt_rd_data_bits_0_9),
    .io_wgt_rd_data_bits_0_10(tensorGemm_io_wgt_rd_data_bits_0_10),
    .io_wgt_rd_data_bits_0_11(tensorGemm_io_wgt_rd_data_bits_0_11),
    .io_wgt_rd_data_bits_0_12(tensorGemm_io_wgt_rd_data_bits_0_12),
    .io_wgt_rd_data_bits_0_13(tensorGemm_io_wgt_rd_data_bits_0_13),
    .io_wgt_rd_data_bits_0_14(tensorGemm_io_wgt_rd_data_bits_0_14),
    .io_wgt_rd_data_bits_0_15(tensorGemm_io_wgt_rd_data_bits_0_15),
    .io_wgt_rd_data_bits_1_0(tensorGemm_io_wgt_rd_data_bits_1_0),
    .io_wgt_rd_data_bits_1_1(tensorGemm_io_wgt_rd_data_bits_1_1),
    .io_wgt_rd_data_bits_1_2(tensorGemm_io_wgt_rd_data_bits_1_2),
    .io_wgt_rd_data_bits_1_3(tensorGemm_io_wgt_rd_data_bits_1_3),
    .io_wgt_rd_data_bits_1_4(tensorGemm_io_wgt_rd_data_bits_1_4),
    .io_wgt_rd_data_bits_1_5(tensorGemm_io_wgt_rd_data_bits_1_5),
    .io_wgt_rd_data_bits_1_6(tensorGemm_io_wgt_rd_data_bits_1_6),
    .io_wgt_rd_data_bits_1_7(tensorGemm_io_wgt_rd_data_bits_1_7),
    .io_wgt_rd_data_bits_1_8(tensorGemm_io_wgt_rd_data_bits_1_8),
    .io_wgt_rd_data_bits_1_9(tensorGemm_io_wgt_rd_data_bits_1_9),
    .io_wgt_rd_data_bits_1_10(tensorGemm_io_wgt_rd_data_bits_1_10),
    .io_wgt_rd_data_bits_1_11(tensorGemm_io_wgt_rd_data_bits_1_11),
    .io_wgt_rd_data_bits_1_12(tensorGemm_io_wgt_rd_data_bits_1_12),
    .io_wgt_rd_data_bits_1_13(tensorGemm_io_wgt_rd_data_bits_1_13),
    .io_wgt_rd_data_bits_1_14(tensorGemm_io_wgt_rd_data_bits_1_14),
    .io_wgt_rd_data_bits_1_15(tensorGemm_io_wgt_rd_data_bits_1_15),
    .io_wgt_rd_data_bits_2_0(tensorGemm_io_wgt_rd_data_bits_2_0),
    .io_wgt_rd_data_bits_2_1(tensorGemm_io_wgt_rd_data_bits_2_1),
    .io_wgt_rd_data_bits_2_2(tensorGemm_io_wgt_rd_data_bits_2_2),
    .io_wgt_rd_data_bits_2_3(tensorGemm_io_wgt_rd_data_bits_2_3),
    .io_wgt_rd_data_bits_2_4(tensorGemm_io_wgt_rd_data_bits_2_4),
    .io_wgt_rd_data_bits_2_5(tensorGemm_io_wgt_rd_data_bits_2_5),
    .io_wgt_rd_data_bits_2_6(tensorGemm_io_wgt_rd_data_bits_2_6),
    .io_wgt_rd_data_bits_2_7(tensorGemm_io_wgt_rd_data_bits_2_7),
    .io_wgt_rd_data_bits_2_8(tensorGemm_io_wgt_rd_data_bits_2_8),
    .io_wgt_rd_data_bits_2_9(tensorGemm_io_wgt_rd_data_bits_2_9),
    .io_wgt_rd_data_bits_2_10(tensorGemm_io_wgt_rd_data_bits_2_10),
    .io_wgt_rd_data_bits_2_11(tensorGemm_io_wgt_rd_data_bits_2_11),
    .io_wgt_rd_data_bits_2_12(tensorGemm_io_wgt_rd_data_bits_2_12),
    .io_wgt_rd_data_bits_2_13(tensorGemm_io_wgt_rd_data_bits_2_13),
    .io_wgt_rd_data_bits_2_14(tensorGemm_io_wgt_rd_data_bits_2_14),
    .io_wgt_rd_data_bits_2_15(tensorGemm_io_wgt_rd_data_bits_2_15),
    .io_wgt_rd_data_bits_3_0(tensorGemm_io_wgt_rd_data_bits_3_0),
    .io_wgt_rd_data_bits_3_1(tensorGemm_io_wgt_rd_data_bits_3_1),
    .io_wgt_rd_data_bits_3_2(tensorGemm_io_wgt_rd_data_bits_3_2),
    .io_wgt_rd_data_bits_3_3(tensorGemm_io_wgt_rd_data_bits_3_3),
    .io_wgt_rd_data_bits_3_4(tensorGemm_io_wgt_rd_data_bits_3_4),
    .io_wgt_rd_data_bits_3_5(tensorGemm_io_wgt_rd_data_bits_3_5),
    .io_wgt_rd_data_bits_3_6(tensorGemm_io_wgt_rd_data_bits_3_6),
    .io_wgt_rd_data_bits_3_7(tensorGemm_io_wgt_rd_data_bits_3_7),
    .io_wgt_rd_data_bits_3_8(tensorGemm_io_wgt_rd_data_bits_3_8),
    .io_wgt_rd_data_bits_3_9(tensorGemm_io_wgt_rd_data_bits_3_9),
    .io_wgt_rd_data_bits_3_10(tensorGemm_io_wgt_rd_data_bits_3_10),
    .io_wgt_rd_data_bits_3_11(tensorGemm_io_wgt_rd_data_bits_3_11),
    .io_wgt_rd_data_bits_3_12(tensorGemm_io_wgt_rd_data_bits_3_12),
    .io_wgt_rd_data_bits_3_13(tensorGemm_io_wgt_rd_data_bits_3_13),
    .io_wgt_rd_data_bits_3_14(tensorGemm_io_wgt_rd_data_bits_3_14),
    .io_wgt_rd_data_bits_3_15(tensorGemm_io_wgt_rd_data_bits_3_15),
    .io_wgt_rd_data_bits_4_0(tensorGemm_io_wgt_rd_data_bits_4_0),
    .io_wgt_rd_data_bits_4_1(tensorGemm_io_wgt_rd_data_bits_4_1),
    .io_wgt_rd_data_bits_4_2(tensorGemm_io_wgt_rd_data_bits_4_2),
    .io_wgt_rd_data_bits_4_3(tensorGemm_io_wgt_rd_data_bits_4_3),
    .io_wgt_rd_data_bits_4_4(tensorGemm_io_wgt_rd_data_bits_4_4),
    .io_wgt_rd_data_bits_4_5(tensorGemm_io_wgt_rd_data_bits_4_5),
    .io_wgt_rd_data_bits_4_6(tensorGemm_io_wgt_rd_data_bits_4_6),
    .io_wgt_rd_data_bits_4_7(tensorGemm_io_wgt_rd_data_bits_4_7),
    .io_wgt_rd_data_bits_4_8(tensorGemm_io_wgt_rd_data_bits_4_8),
    .io_wgt_rd_data_bits_4_9(tensorGemm_io_wgt_rd_data_bits_4_9),
    .io_wgt_rd_data_bits_4_10(tensorGemm_io_wgt_rd_data_bits_4_10),
    .io_wgt_rd_data_bits_4_11(tensorGemm_io_wgt_rd_data_bits_4_11),
    .io_wgt_rd_data_bits_4_12(tensorGemm_io_wgt_rd_data_bits_4_12),
    .io_wgt_rd_data_bits_4_13(tensorGemm_io_wgt_rd_data_bits_4_13),
    .io_wgt_rd_data_bits_4_14(tensorGemm_io_wgt_rd_data_bits_4_14),
    .io_wgt_rd_data_bits_4_15(tensorGemm_io_wgt_rd_data_bits_4_15),
    .io_wgt_rd_data_bits_5_0(tensorGemm_io_wgt_rd_data_bits_5_0),
    .io_wgt_rd_data_bits_5_1(tensorGemm_io_wgt_rd_data_bits_5_1),
    .io_wgt_rd_data_bits_5_2(tensorGemm_io_wgt_rd_data_bits_5_2),
    .io_wgt_rd_data_bits_5_3(tensorGemm_io_wgt_rd_data_bits_5_3),
    .io_wgt_rd_data_bits_5_4(tensorGemm_io_wgt_rd_data_bits_5_4),
    .io_wgt_rd_data_bits_5_5(tensorGemm_io_wgt_rd_data_bits_5_5),
    .io_wgt_rd_data_bits_5_6(tensorGemm_io_wgt_rd_data_bits_5_6),
    .io_wgt_rd_data_bits_5_7(tensorGemm_io_wgt_rd_data_bits_5_7),
    .io_wgt_rd_data_bits_5_8(tensorGemm_io_wgt_rd_data_bits_5_8),
    .io_wgt_rd_data_bits_5_9(tensorGemm_io_wgt_rd_data_bits_5_9),
    .io_wgt_rd_data_bits_5_10(tensorGemm_io_wgt_rd_data_bits_5_10),
    .io_wgt_rd_data_bits_5_11(tensorGemm_io_wgt_rd_data_bits_5_11),
    .io_wgt_rd_data_bits_5_12(tensorGemm_io_wgt_rd_data_bits_5_12),
    .io_wgt_rd_data_bits_5_13(tensorGemm_io_wgt_rd_data_bits_5_13),
    .io_wgt_rd_data_bits_5_14(tensorGemm_io_wgt_rd_data_bits_5_14),
    .io_wgt_rd_data_bits_5_15(tensorGemm_io_wgt_rd_data_bits_5_15),
    .io_wgt_rd_data_bits_6_0(tensorGemm_io_wgt_rd_data_bits_6_0),
    .io_wgt_rd_data_bits_6_1(tensorGemm_io_wgt_rd_data_bits_6_1),
    .io_wgt_rd_data_bits_6_2(tensorGemm_io_wgt_rd_data_bits_6_2),
    .io_wgt_rd_data_bits_6_3(tensorGemm_io_wgt_rd_data_bits_6_3),
    .io_wgt_rd_data_bits_6_4(tensorGemm_io_wgt_rd_data_bits_6_4),
    .io_wgt_rd_data_bits_6_5(tensorGemm_io_wgt_rd_data_bits_6_5),
    .io_wgt_rd_data_bits_6_6(tensorGemm_io_wgt_rd_data_bits_6_6),
    .io_wgt_rd_data_bits_6_7(tensorGemm_io_wgt_rd_data_bits_6_7),
    .io_wgt_rd_data_bits_6_8(tensorGemm_io_wgt_rd_data_bits_6_8),
    .io_wgt_rd_data_bits_6_9(tensorGemm_io_wgt_rd_data_bits_6_9),
    .io_wgt_rd_data_bits_6_10(tensorGemm_io_wgt_rd_data_bits_6_10),
    .io_wgt_rd_data_bits_6_11(tensorGemm_io_wgt_rd_data_bits_6_11),
    .io_wgt_rd_data_bits_6_12(tensorGemm_io_wgt_rd_data_bits_6_12),
    .io_wgt_rd_data_bits_6_13(tensorGemm_io_wgt_rd_data_bits_6_13),
    .io_wgt_rd_data_bits_6_14(tensorGemm_io_wgt_rd_data_bits_6_14),
    .io_wgt_rd_data_bits_6_15(tensorGemm_io_wgt_rd_data_bits_6_15),
    .io_wgt_rd_data_bits_7_0(tensorGemm_io_wgt_rd_data_bits_7_0),
    .io_wgt_rd_data_bits_7_1(tensorGemm_io_wgt_rd_data_bits_7_1),
    .io_wgt_rd_data_bits_7_2(tensorGemm_io_wgt_rd_data_bits_7_2),
    .io_wgt_rd_data_bits_7_3(tensorGemm_io_wgt_rd_data_bits_7_3),
    .io_wgt_rd_data_bits_7_4(tensorGemm_io_wgt_rd_data_bits_7_4),
    .io_wgt_rd_data_bits_7_5(tensorGemm_io_wgt_rd_data_bits_7_5),
    .io_wgt_rd_data_bits_7_6(tensorGemm_io_wgt_rd_data_bits_7_6),
    .io_wgt_rd_data_bits_7_7(tensorGemm_io_wgt_rd_data_bits_7_7),
    .io_wgt_rd_data_bits_7_8(tensorGemm_io_wgt_rd_data_bits_7_8),
    .io_wgt_rd_data_bits_7_9(tensorGemm_io_wgt_rd_data_bits_7_9),
    .io_wgt_rd_data_bits_7_10(tensorGemm_io_wgt_rd_data_bits_7_10),
    .io_wgt_rd_data_bits_7_11(tensorGemm_io_wgt_rd_data_bits_7_11),
    .io_wgt_rd_data_bits_7_12(tensorGemm_io_wgt_rd_data_bits_7_12),
    .io_wgt_rd_data_bits_7_13(tensorGemm_io_wgt_rd_data_bits_7_13),
    .io_wgt_rd_data_bits_7_14(tensorGemm_io_wgt_rd_data_bits_7_14),
    .io_wgt_rd_data_bits_7_15(tensorGemm_io_wgt_rd_data_bits_7_15),
    .io_wgt_rd_data_bits_8_0(tensorGemm_io_wgt_rd_data_bits_8_0),
    .io_wgt_rd_data_bits_8_1(tensorGemm_io_wgt_rd_data_bits_8_1),
    .io_wgt_rd_data_bits_8_2(tensorGemm_io_wgt_rd_data_bits_8_2),
    .io_wgt_rd_data_bits_8_3(tensorGemm_io_wgt_rd_data_bits_8_3),
    .io_wgt_rd_data_bits_8_4(tensorGemm_io_wgt_rd_data_bits_8_4),
    .io_wgt_rd_data_bits_8_5(tensorGemm_io_wgt_rd_data_bits_8_5),
    .io_wgt_rd_data_bits_8_6(tensorGemm_io_wgt_rd_data_bits_8_6),
    .io_wgt_rd_data_bits_8_7(tensorGemm_io_wgt_rd_data_bits_8_7),
    .io_wgt_rd_data_bits_8_8(tensorGemm_io_wgt_rd_data_bits_8_8),
    .io_wgt_rd_data_bits_8_9(tensorGemm_io_wgt_rd_data_bits_8_9),
    .io_wgt_rd_data_bits_8_10(tensorGemm_io_wgt_rd_data_bits_8_10),
    .io_wgt_rd_data_bits_8_11(tensorGemm_io_wgt_rd_data_bits_8_11),
    .io_wgt_rd_data_bits_8_12(tensorGemm_io_wgt_rd_data_bits_8_12),
    .io_wgt_rd_data_bits_8_13(tensorGemm_io_wgt_rd_data_bits_8_13),
    .io_wgt_rd_data_bits_8_14(tensorGemm_io_wgt_rd_data_bits_8_14),
    .io_wgt_rd_data_bits_8_15(tensorGemm_io_wgt_rd_data_bits_8_15),
    .io_wgt_rd_data_bits_9_0(tensorGemm_io_wgt_rd_data_bits_9_0),
    .io_wgt_rd_data_bits_9_1(tensorGemm_io_wgt_rd_data_bits_9_1),
    .io_wgt_rd_data_bits_9_2(tensorGemm_io_wgt_rd_data_bits_9_2),
    .io_wgt_rd_data_bits_9_3(tensorGemm_io_wgt_rd_data_bits_9_3),
    .io_wgt_rd_data_bits_9_4(tensorGemm_io_wgt_rd_data_bits_9_4),
    .io_wgt_rd_data_bits_9_5(tensorGemm_io_wgt_rd_data_bits_9_5),
    .io_wgt_rd_data_bits_9_6(tensorGemm_io_wgt_rd_data_bits_9_6),
    .io_wgt_rd_data_bits_9_7(tensorGemm_io_wgt_rd_data_bits_9_7),
    .io_wgt_rd_data_bits_9_8(tensorGemm_io_wgt_rd_data_bits_9_8),
    .io_wgt_rd_data_bits_9_9(tensorGemm_io_wgt_rd_data_bits_9_9),
    .io_wgt_rd_data_bits_9_10(tensorGemm_io_wgt_rd_data_bits_9_10),
    .io_wgt_rd_data_bits_9_11(tensorGemm_io_wgt_rd_data_bits_9_11),
    .io_wgt_rd_data_bits_9_12(tensorGemm_io_wgt_rd_data_bits_9_12),
    .io_wgt_rd_data_bits_9_13(tensorGemm_io_wgt_rd_data_bits_9_13),
    .io_wgt_rd_data_bits_9_14(tensorGemm_io_wgt_rd_data_bits_9_14),
    .io_wgt_rd_data_bits_9_15(tensorGemm_io_wgt_rd_data_bits_9_15),
    .io_wgt_rd_data_bits_10_0(tensorGemm_io_wgt_rd_data_bits_10_0),
    .io_wgt_rd_data_bits_10_1(tensorGemm_io_wgt_rd_data_bits_10_1),
    .io_wgt_rd_data_bits_10_2(tensorGemm_io_wgt_rd_data_bits_10_2),
    .io_wgt_rd_data_bits_10_3(tensorGemm_io_wgt_rd_data_bits_10_3),
    .io_wgt_rd_data_bits_10_4(tensorGemm_io_wgt_rd_data_bits_10_4),
    .io_wgt_rd_data_bits_10_5(tensorGemm_io_wgt_rd_data_bits_10_5),
    .io_wgt_rd_data_bits_10_6(tensorGemm_io_wgt_rd_data_bits_10_6),
    .io_wgt_rd_data_bits_10_7(tensorGemm_io_wgt_rd_data_bits_10_7),
    .io_wgt_rd_data_bits_10_8(tensorGemm_io_wgt_rd_data_bits_10_8),
    .io_wgt_rd_data_bits_10_9(tensorGemm_io_wgt_rd_data_bits_10_9),
    .io_wgt_rd_data_bits_10_10(tensorGemm_io_wgt_rd_data_bits_10_10),
    .io_wgt_rd_data_bits_10_11(tensorGemm_io_wgt_rd_data_bits_10_11),
    .io_wgt_rd_data_bits_10_12(tensorGemm_io_wgt_rd_data_bits_10_12),
    .io_wgt_rd_data_bits_10_13(tensorGemm_io_wgt_rd_data_bits_10_13),
    .io_wgt_rd_data_bits_10_14(tensorGemm_io_wgt_rd_data_bits_10_14),
    .io_wgt_rd_data_bits_10_15(tensorGemm_io_wgt_rd_data_bits_10_15),
    .io_wgt_rd_data_bits_11_0(tensorGemm_io_wgt_rd_data_bits_11_0),
    .io_wgt_rd_data_bits_11_1(tensorGemm_io_wgt_rd_data_bits_11_1),
    .io_wgt_rd_data_bits_11_2(tensorGemm_io_wgt_rd_data_bits_11_2),
    .io_wgt_rd_data_bits_11_3(tensorGemm_io_wgt_rd_data_bits_11_3),
    .io_wgt_rd_data_bits_11_4(tensorGemm_io_wgt_rd_data_bits_11_4),
    .io_wgt_rd_data_bits_11_5(tensorGemm_io_wgt_rd_data_bits_11_5),
    .io_wgt_rd_data_bits_11_6(tensorGemm_io_wgt_rd_data_bits_11_6),
    .io_wgt_rd_data_bits_11_7(tensorGemm_io_wgt_rd_data_bits_11_7),
    .io_wgt_rd_data_bits_11_8(tensorGemm_io_wgt_rd_data_bits_11_8),
    .io_wgt_rd_data_bits_11_9(tensorGemm_io_wgt_rd_data_bits_11_9),
    .io_wgt_rd_data_bits_11_10(tensorGemm_io_wgt_rd_data_bits_11_10),
    .io_wgt_rd_data_bits_11_11(tensorGemm_io_wgt_rd_data_bits_11_11),
    .io_wgt_rd_data_bits_11_12(tensorGemm_io_wgt_rd_data_bits_11_12),
    .io_wgt_rd_data_bits_11_13(tensorGemm_io_wgt_rd_data_bits_11_13),
    .io_wgt_rd_data_bits_11_14(tensorGemm_io_wgt_rd_data_bits_11_14),
    .io_wgt_rd_data_bits_11_15(tensorGemm_io_wgt_rd_data_bits_11_15),
    .io_wgt_rd_data_bits_12_0(tensorGemm_io_wgt_rd_data_bits_12_0),
    .io_wgt_rd_data_bits_12_1(tensorGemm_io_wgt_rd_data_bits_12_1),
    .io_wgt_rd_data_bits_12_2(tensorGemm_io_wgt_rd_data_bits_12_2),
    .io_wgt_rd_data_bits_12_3(tensorGemm_io_wgt_rd_data_bits_12_3),
    .io_wgt_rd_data_bits_12_4(tensorGemm_io_wgt_rd_data_bits_12_4),
    .io_wgt_rd_data_bits_12_5(tensorGemm_io_wgt_rd_data_bits_12_5),
    .io_wgt_rd_data_bits_12_6(tensorGemm_io_wgt_rd_data_bits_12_6),
    .io_wgt_rd_data_bits_12_7(tensorGemm_io_wgt_rd_data_bits_12_7),
    .io_wgt_rd_data_bits_12_8(tensorGemm_io_wgt_rd_data_bits_12_8),
    .io_wgt_rd_data_bits_12_9(tensorGemm_io_wgt_rd_data_bits_12_9),
    .io_wgt_rd_data_bits_12_10(tensorGemm_io_wgt_rd_data_bits_12_10),
    .io_wgt_rd_data_bits_12_11(tensorGemm_io_wgt_rd_data_bits_12_11),
    .io_wgt_rd_data_bits_12_12(tensorGemm_io_wgt_rd_data_bits_12_12),
    .io_wgt_rd_data_bits_12_13(tensorGemm_io_wgt_rd_data_bits_12_13),
    .io_wgt_rd_data_bits_12_14(tensorGemm_io_wgt_rd_data_bits_12_14),
    .io_wgt_rd_data_bits_12_15(tensorGemm_io_wgt_rd_data_bits_12_15),
    .io_wgt_rd_data_bits_13_0(tensorGemm_io_wgt_rd_data_bits_13_0),
    .io_wgt_rd_data_bits_13_1(tensorGemm_io_wgt_rd_data_bits_13_1),
    .io_wgt_rd_data_bits_13_2(tensorGemm_io_wgt_rd_data_bits_13_2),
    .io_wgt_rd_data_bits_13_3(tensorGemm_io_wgt_rd_data_bits_13_3),
    .io_wgt_rd_data_bits_13_4(tensorGemm_io_wgt_rd_data_bits_13_4),
    .io_wgt_rd_data_bits_13_5(tensorGemm_io_wgt_rd_data_bits_13_5),
    .io_wgt_rd_data_bits_13_6(tensorGemm_io_wgt_rd_data_bits_13_6),
    .io_wgt_rd_data_bits_13_7(tensorGemm_io_wgt_rd_data_bits_13_7),
    .io_wgt_rd_data_bits_13_8(tensorGemm_io_wgt_rd_data_bits_13_8),
    .io_wgt_rd_data_bits_13_9(tensorGemm_io_wgt_rd_data_bits_13_9),
    .io_wgt_rd_data_bits_13_10(tensorGemm_io_wgt_rd_data_bits_13_10),
    .io_wgt_rd_data_bits_13_11(tensorGemm_io_wgt_rd_data_bits_13_11),
    .io_wgt_rd_data_bits_13_12(tensorGemm_io_wgt_rd_data_bits_13_12),
    .io_wgt_rd_data_bits_13_13(tensorGemm_io_wgt_rd_data_bits_13_13),
    .io_wgt_rd_data_bits_13_14(tensorGemm_io_wgt_rd_data_bits_13_14),
    .io_wgt_rd_data_bits_13_15(tensorGemm_io_wgt_rd_data_bits_13_15),
    .io_wgt_rd_data_bits_14_0(tensorGemm_io_wgt_rd_data_bits_14_0),
    .io_wgt_rd_data_bits_14_1(tensorGemm_io_wgt_rd_data_bits_14_1),
    .io_wgt_rd_data_bits_14_2(tensorGemm_io_wgt_rd_data_bits_14_2),
    .io_wgt_rd_data_bits_14_3(tensorGemm_io_wgt_rd_data_bits_14_3),
    .io_wgt_rd_data_bits_14_4(tensorGemm_io_wgt_rd_data_bits_14_4),
    .io_wgt_rd_data_bits_14_5(tensorGemm_io_wgt_rd_data_bits_14_5),
    .io_wgt_rd_data_bits_14_6(tensorGemm_io_wgt_rd_data_bits_14_6),
    .io_wgt_rd_data_bits_14_7(tensorGemm_io_wgt_rd_data_bits_14_7),
    .io_wgt_rd_data_bits_14_8(tensorGemm_io_wgt_rd_data_bits_14_8),
    .io_wgt_rd_data_bits_14_9(tensorGemm_io_wgt_rd_data_bits_14_9),
    .io_wgt_rd_data_bits_14_10(tensorGemm_io_wgt_rd_data_bits_14_10),
    .io_wgt_rd_data_bits_14_11(tensorGemm_io_wgt_rd_data_bits_14_11),
    .io_wgt_rd_data_bits_14_12(tensorGemm_io_wgt_rd_data_bits_14_12),
    .io_wgt_rd_data_bits_14_13(tensorGemm_io_wgt_rd_data_bits_14_13),
    .io_wgt_rd_data_bits_14_14(tensorGemm_io_wgt_rd_data_bits_14_14),
    .io_wgt_rd_data_bits_14_15(tensorGemm_io_wgt_rd_data_bits_14_15),
    .io_wgt_rd_data_bits_15_0(tensorGemm_io_wgt_rd_data_bits_15_0),
    .io_wgt_rd_data_bits_15_1(tensorGemm_io_wgt_rd_data_bits_15_1),
    .io_wgt_rd_data_bits_15_2(tensorGemm_io_wgt_rd_data_bits_15_2),
    .io_wgt_rd_data_bits_15_3(tensorGemm_io_wgt_rd_data_bits_15_3),
    .io_wgt_rd_data_bits_15_4(tensorGemm_io_wgt_rd_data_bits_15_4),
    .io_wgt_rd_data_bits_15_5(tensorGemm_io_wgt_rd_data_bits_15_5),
    .io_wgt_rd_data_bits_15_6(tensorGemm_io_wgt_rd_data_bits_15_6),
    .io_wgt_rd_data_bits_15_7(tensorGemm_io_wgt_rd_data_bits_15_7),
    .io_wgt_rd_data_bits_15_8(tensorGemm_io_wgt_rd_data_bits_15_8),
    .io_wgt_rd_data_bits_15_9(tensorGemm_io_wgt_rd_data_bits_15_9),
    .io_wgt_rd_data_bits_15_10(tensorGemm_io_wgt_rd_data_bits_15_10),
    .io_wgt_rd_data_bits_15_11(tensorGemm_io_wgt_rd_data_bits_15_11),
    .io_wgt_rd_data_bits_15_12(tensorGemm_io_wgt_rd_data_bits_15_12),
    .io_wgt_rd_data_bits_15_13(tensorGemm_io_wgt_rd_data_bits_15_13),
    .io_wgt_rd_data_bits_15_14(tensorGemm_io_wgt_rd_data_bits_15_14),
    .io_wgt_rd_data_bits_15_15(tensorGemm_io_wgt_rd_data_bits_15_15),
    .io_acc_rd_idx_valid(tensorGemm_io_acc_rd_idx_valid),
    .io_acc_rd_idx_bits(tensorGemm_io_acc_rd_idx_bits),
    .io_acc_rd_data_valid(tensorGemm_io_acc_rd_data_valid),
    .io_acc_rd_data_bits_0_0(tensorGemm_io_acc_rd_data_bits_0_0),
    .io_acc_rd_data_bits_0_1(tensorGemm_io_acc_rd_data_bits_0_1),
    .io_acc_rd_data_bits_0_2(tensorGemm_io_acc_rd_data_bits_0_2),
    .io_acc_rd_data_bits_0_3(tensorGemm_io_acc_rd_data_bits_0_3),
    .io_acc_rd_data_bits_0_4(tensorGemm_io_acc_rd_data_bits_0_4),
    .io_acc_rd_data_bits_0_5(tensorGemm_io_acc_rd_data_bits_0_5),
    .io_acc_rd_data_bits_0_6(tensorGemm_io_acc_rd_data_bits_0_6),
    .io_acc_rd_data_bits_0_7(tensorGemm_io_acc_rd_data_bits_0_7),
    .io_acc_rd_data_bits_0_8(tensorGemm_io_acc_rd_data_bits_0_8),
    .io_acc_rd_data_bits_0_9(tensorGemm_io_acc_rd_data_bits_0_9),
    .io_acc_rd_data_bits_0_10(tensorGemm_io_acc_rd_data_bits_0_10),
    .io_acc_rd_data_bits_0_11(tensorGemm_io_acc_rd_data_bits_0_11),
    .io_acc_rd_data_bits_0_12(tensorGemm_io_acc_rd_data_bits_0_12),
    .io_acc_rd_data_bits_0_13(tensorGemm_io_acc_rd_data_bits_0_13),
    .io_acc_rd_data_bits_0_14(tensorGemm_io_acc_rd_data_bits_0_14),
    .io_acc_rd_data_bits_0_15(tensorGemm_io_acc_rd_data_bits_0_15),
    .io_acc_wr_valid(tensorGemm_io_acc_wr_valid),
    .io_acc_wr_bits_idx(tensorGemm_io_acc_wr_bits_idx),
    .io_acc_wr_bits_data_0_0(tensorGemm_io_acc_wr_bits_data_0_0),
    .io_acc_wr_bits_data_0_1(tensorGemm_io_acc_wr_bits_data_0_1),
    .io_acc_wr_bits_data_0_2(tensorGemm_io_acc_wr_bits_data_0_2),
    .io_acc_wr_bits_data_0_3(tensorGemm_io_acc_wr_bits_data_0_3),
    .io_acc_wr_bits_data_0_4(tensorGemm_io_acc_wr_bits_data_0_4),
    .io_acc_wr_bits_data_0_5(tensorGemm_io_acc_wr_bits_data_0_5),
    .io_acc_wr_bits_data_0_6(tensorGemm_io_acc_wr_bits_data_0_6),
    .io_acc_wr_bits_data_0_7(tensorGemm_io_acc_wr_bits_data_0_7),
    .io_acc_wr_bits_data_0_8(tensorGemm_io_acc_wr_bits_data_0_8),
    .io_acc_wr_bits_data_0_9(tensorGemm_io_acc_wr_bits_data_0_9),
    .io_acc_wr_bits_data_0_10(tensorGemm_io_acc_wr_bits_data_0_10),
    .io_acc_wr_bits_data_0_11(tensorGemm_io_acc_wr_bits_data_0_11),
    .io_acc_wr_bits_data_0_12(tensorGemm_io_acc_wr_bits_data_0_12),
    .io_acc_wr_bits_data_0_13(tensorGemm_io_acc_wr_bits_data_0_13),
    .io_acc_wr_bits_data_0_14(tensorGemm_io_acc_wr_bits_data_0_14),
    .io_acc_wr_bits_data_0_15(tensorGemm_io_acc_wr_bits_data_0_15),
    .io_out_wr_valid(tensorGemm_io_out_wr_valid),
    .io_out_wr_bits_idx(tensorGemm_io_out_wr_bits_idx),
    .io_out_wr_bits_data_0_0(tensorGemm_io_out_wr_bits_data_0_0),
    .io_out_wr_bits_data_0_1(tensorGemm_io_out_wr_bits_data_0_1),
    .io_out_wr_bits_data_0_2(tensorGemm_io_out_wr_bits_data_0_2),
    .io_out_wr_bits_data_0_3(tensorGemm_io_out_wr_bits_data_0_3),
    .io_out_wr_bits_data_0_4(tensorGemm_io_out_wr_bits_data_0_4),
    .io_out_wr_bits_data_0_5(tensorGemm_io_out_wr_bits_data_0_5),
    .io_out_wr_bits_data_0_6(tensorGemm_io_out_wr_bits_data_0_6),
    .io_out_wr_bits_data_0_7(tensorGemm_io_out_wr_bits_data_0_7),
    .io_out_wr_bits_data_0_8(tensorGemm_io_out_wr_bits_data_0_8),
    .io_out_wr_bits_data_0_9(tensorGemm_io_out_wr_bits_data_0_9),
    .io_out_wr_bits_data_0_10(tensorGemm_io_out_wr_bits_data_0_10),
    .io_out_wr_bits_data_0_11(tensorGemm_io_out_wr_bits_data_0_11),
    .io_out_wr_bits_data_0_12(tensorGemm_io_out_wr_bits_data_0_12),
    .io_out_wr_bits_data_0_13(tensorGemm_io_out_wr_bits_data_0_13),
    .io_out_wr_bits_data_0_14(tensorGemm_io_out_wr_bits_data_0_14),
    .io_out_wr_bits_data_0_15(tensorGemm_io_out_wr_bits_data_0_15)
  );
  TensorAlu tensorAlu ( // @[Compute.scala 59:25:@22768.4]
    .clock(tensorAlu_clock),
    .reset(tensorAlu_reset),
    .io_start(tensorAlu_io_start),
    .io_done(tensorAlu_io_done),
    .io_inst(tensorAlu_io_inst),
    .io_uop_idx_valid(tensorAlu_io_uop_idx_valid),
    .io_uop_idx_bits(tensorAlu_io_uop_idx_bits),
    .io_uop_data_valid(tensorAlu_io_uop_data_valid),
    .io_uop_data_bits_u1(tensorAlu_io_uop_data_bits_u1),
    .io_uop_data_bits_u0(tensorAlu_io_uop_data_bits_u0),
    .io_acc_rd_idx_valid(tensorAlu_io_acc_rd_idx_valid),
    .io_acc_rd_idx_bits(tensorAlu_io_acc_rd_idx_bits),
    .io_acc_rd_data_valid(tensorAlu_io_acc_rd_data_valid),
    .io_acc_rd_data_bits_0_0(tensorAlu_io_acc_rd_data_bits_0_0),
    .io_acc_rd_data_bits_0_1(tensorAlu_io_acc_rd_data_bits_0_1),
    .io_acc_rd_data_bits_0_2(tensorAlu_io_acc_rd_data_bits_0_2),
    .io_acc_rd_data_bits_0_3(tensorAlu_io_acc_rd_data_bits_0_3),
    .io_acc_rd_data_bits_0_4(tensorAlu_io_acc_rd_data_bits_0_4),
    .io_acc_rd_data_bits_0_5(tensorAlu_io_acc_rd_data_bits_0_5),
    .io_acc_rd_data_bits_0_6(tensorAlu_io_acc_rd_data_bits_0_6),
    .io_acc_rd_data_bits_0_7(tensorAlu_io_acc_rd_data_bits_0_7),
    .io_acc_rd_data_bits_0_8(tensorAlu_io_acc_rd_data_bits_0_8),
    .io_acc_rd_data_bits_0_9(tensorAlu_io_acc_rd_data_bits_0_9),
    .io_acc_rd_data_bits_0_10(tensorAlu_io_acc_rd_data_bits_0_10),
    .io_acc_rd_data_bits_0_11(tensorAlu_io_acc_rd_data_bits_0_11),
    .io_acc_rd_data_bits_0_12(tensorAlu_io_acc_rd_data_bits_0_12),
    .io_acc_rd_data_bits_0_13(tensorAlu_io_acc_rd_data_bits_0_13),
    .io_acc_rd_data_bits_0_14(tensorAlu_io_acc_rd_data_bits_0_14),
    .io_acc_rd_data_bits_0_15(tensorAlu_io_acc_rd_data_bits_0_15),
    .io_acc_wr_valid(tensorAlu_io_acc_wr_valid),
    .io_acc_wr_bits_idx(tensorAlu_io_acc_wr_bits_idx),
    .io_acc_wr_bits_data_0_0(tensorAlu_io_acc_wr_bits_data_0_0),
    .io_acc_wr_bits_data_0_1(tensorAlu_io_acc_wr_bits_data_0_1),
    .io_acc_wr_bits_data_0_2(tensorAlu_io_acc_wr_bits_data_0_2),
    .io_acc_wr_bits_data_0_3(tensorAlu_io_acc_wr_bits_data_0_3),
    .io_acc_wr_bits_data_0_4(tensorAlu_io_acc_wr_bits_data_0_4),
    .io_acc_wr_bits_data_0_5(tensorAlu_io_acc_wr_bits_data_0_5),
    .io_acc_wr_bits_data_0_6(tensorAlu_io_acc_wr_bits_data_0_6),
    .io_acc_wr_bits_data_0_7(tensorAlu_io_acc_wr_bits_data_0_7),
    .io_acc_wr_bits_data_0_8(tensorAlu_io_acc_wr_bits_data_0_8),
    .io_acc_wr_bits_data_0_9(tensorAlu_io_acc_wr_bits_data_0_9),
    .io_acc_wr_bits_data_0_10(tensorAlu_io_acc_wr_bits_data_0_10),
    .io_acc_wr_bits_data_0_11(tensorAlu_io_acc_wr_bits_data_0_11),
    .io_acc_wr_bits_data_0_12(tensorAlu_io_acc_wr_bits_data_0_12),
    .io_acc_wr_bits_data_0_13(tensorAlu_io_acc_wr_bits_data_0_13),
    .io_acc_wr_bits_data_0_14(tensorAlu_io_acc_wr_bits_data_0_14),
    .io_acc_wr_bits_data_0_15(tensorAlu_io_acc_wr_bits_data_0_15),
    .io_out_wr_valid(tensorAlu_io_out_wr_valid),
    .io_out_wr_bits_idx(tensorAlu_io_out_wr_bits_idx),
    .io_out_wr_bits_data_0_0(tensorAlu_io_out_wr_bits_data_0_0),
    .io_out_wr_bits_data_0_1(tensorAlu_io_out_wr_bits_data_0_1),
    .io_out_wr_bits_data_0_2(tensorAlu_io_out_wr_bits_data_0_2),
    .io_out_wr_bits_data_0_3(tensorAlu_io_out_wr_bits_data_0_3),
    .io_out_wr_bits_data_0_4(tensorAlu_io_out_wr_bits_data_0_4),
    .io_out_wr_bits_data_0_5(tensorAlu_io_out_wr_bits_data_0_5),
    .io_out_wr_bits_data_0_6(tensorAlu_io_out_wr_bits_data_0_6),
    .io_out_wr_bits_data_0_7(tensorAlu_io_out_wr_bits_data_0_7),
    .io_out_wr_bits_data_0_8(tensorAlu_io_out_wr_bits_data_0_8),
    .io_out_wr_bits_data_0_9(tensorAlu_io_out_wr_bits_data_0_9),
    .io_out_wr_bits_data_0_10(tensorAlu_io_out_wr_bits_data_0_10),
    .io_out_wr_bits_data_0_11(tensorAlu_io_out_wr_bits_data_0_11),
    .io_out_wr_bits_data_0_12(tensorAlu_io_out_wr_bits_data_0_12),
    .io_out_wr_bits_data_0_13(tensorAlu_io_out_wr_bits_data_0_13),
    .io_out_wr_bits_data_0_14(tensorAlu_io_out_wr_bits_data_0_14),
    .io_out_wr_bits_data_0_15(tensorAlu_io_out_wr_bits_data_0_15)
  );
  Queue_1 inst_q ( // @[Compute.scala 61:22:@22771.4]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits)
  );
  ComputeDecode dec ( // @[Compute.scala 64:19:@22774.4]
    .io_inst(dec_io_inst),
    .io_push_next(dec_io_push_next),
    .io_push_prev(dec_io_push_prev),
    .io_pop_next(dec_io_pop_next),
    .io_pop_prev(dec_io_pop_prev),
    .io_isLoadAcc(dec_io_isLoadAcc),
    .io_isLoadUop(dec_io_isLoadUop),
    .io_isSync(dec_io_isSync),
    .io_isAlu(dec_io_isAlu),
    .io_isGemm(dec_io_isGemm),
    .io_isFinish(dec_io_isFinish)
  );
  assign inst_type = {dec_io_isFinish,dec_io_isAlu,dec_io_isGemm,dec_io_isLoadAcc,dec_io_isLoadUop}; // @[Cat.scala 30:58:@22781.4]
  assign _T_7054 = dec_io_pop_prev ? s_0_io_sready : 1'h1; // @[Compute.scala 74:40:@22782.4]
  assign sprev = inst_q_io_deq_valid & _T_7054; // @[Compute.scala 74:35:@22783.4]
  assign _T_7056 = dec_io_pop_next ? s_1_io_sready : 1'h1; // @[Compute.scala 75:40:@22784.4]
  assign snext = inst_q_io_deq_valid & _T_7056; // @[Compute.scala 75:35:@22785.4]
  assign start = snext & sprev; // @[Compute.scala 76:21:@22786.4]
  assign _T_7064 = 5'h10 == inst_type; // @[Mux.scala 46:19:@22787.4]
  assign _T_7066 = 5'h8 == inst_type; // @[Mux.scala 46:19:@22789.4]
  assign _T_7067 = _T_7066 ? tensorAlu_io_done : _T_7064; // @[Mux.scala 46:16:@22790.4]
  assign _T_7068 = 5'h4 == inst_type; // @[Mux.scala 46:19:@22791.4]
  assign _T_7069 = _T_7068 ? tensorGemm_io_done : _T_7067; // @[Mux.scala 46:16:@22792.4]
  assign _T_7070 = 5'h2 == inst_type; // @[Mux.scala 46:19:@22793.4]
  assign _T_7071 = _T_7070 ? tensorAcc_io_done : _T_7069; // @[Mux.scala 46:16:@22794.4]
  assign _T_7072 = 5'h1 == inst_type; // @[Mux.scala 46:19:@22795.4]
  assign done = _T_7072 ? loadUop_io_done : _T_7071; // @[Mux.scala 46:16:@22796.4]
  assign _T_7073 = 2'h0 == state; // @[Conditional.scala 37:30:@22797.4]
  assign _T_7075 = inst_type != 5'h0; // @[Compute.scala 96:30:@22804.10]
  assign _GEN_0 = _T_7075 ? 2'h2 : state; // @[Compute.scala 96:35:@22805.10]
  assign _GEN_1 = dec_io_isSync ? 2'h1 : _GEN_0; // @[Compute.scala 94:29:@22800.8]
  assign _GEN_2 = start ? _GEN_1 : state; // @[Compute.scala 93:19:@22799.6]
  assign _T_7076 = 2'h1 == state; // @[Conditional.scala 37:30:@22811.6]
  assign _T_7077 = 2'h2 == state; // @[Conditional.scala 37:30:@22816.8]
  assign _GEN_3 = done ? 2'h0 : state; // @[Compute.scala 105:18:@22818.10]
  assign _GEN_4 = _T_7077 ? _GEN_3 : state; // @[Conditional.scala 39:67:@22817.8]
  assign _GEN_5 = _T_7076 ? 2'h0 : _GEN_4; // @[Conditional.scala 39:67:@22812.6]
  assign _GEN_6 = _T_7073 ? _GEN_2 : _GEN_5; // @[Conditional.scala 40:58:@22798.4]
  assign _T_7078 = state == 2'h2; // @[Compute.scala 113:33:@22825.4]
  assign _T_7079 = _T_7078 & done; // @[Compute.scala 113:42:@22826.4]
  assign _T_7080 = state == 2'h1; // @[Compute.scala 113:59:@22827.4]
  assign _T_7081 = _T_7079 | _T_7080; // @[Compute.scala 113:50:@22828.4]
  assign _T_7082 = state == 2'h0; // @[Compute.scala 116:29:@22830.4]
  assign _T_7083 = _T_7082 & start; // @[Compute.scala 116:39:@22831.4]
  assign io_o_post_0 = dec_io_push_prev & _T_7081; // @[Compute.scala 164:16:@23565.4]
  assign io_o_post_1 = dec_io_push_next & _T_7081; // @[Compute.scala 165:16:@23571.4]
  assign io_inst_ready = inst_q_io_enq_ready; // @[Compute.scala 112:17:@22824.4]
  assign io_vme_rd_0_cmd_valid = loadUop_io_vme_rd_cmd_valid; // @[Compute.scala 119:16:@22841.4]
  assign io_vme_rd_0_cmd_bits_addr = loadUop_io_vme_rd_cmd_bits_addr; // @[Compute.scala 119:16:@22840.4]
  assign io_vme_rd_0_cmd_bits_len = loadUop_io_vme_rd_cmd_bits_len; // @[Compute.scala 119:16:@22839.4]
  assign io_vme_rd_0_data_ready = loadUop_io_vme_rd_data_ready; // @[Compute.scala 119:16:@22838.4]
  assign io_vme_rd_1_cmd_valid = tensorAcc_io_vme_rd_cmd_valid; // @[Compute.scala 128:16:@22879.4]
  assign io_vme_rd_1_cmd_bits_addr = tensorAcc_io_vme_rd_cmd_bits_addr; // @[Compute.scala 128:16:@22878.4]
  assign io_vme_rd_1_cmd_bits_len = tensorAcc_io_vme_rd_cmd_bits_len; // @[Compute.scala 128:16:@22877.4]
  assign io_vme_rd_1_data_ready = tensorAcc_io_vme_rd_data_ready; // @[Compute.scala 128:16:@22876.4]
  assign io_inp_rd_idx_valid = tensorGemm_io_inp_rd_idx_valid; // @[Compute.scala 136:21:@22928.4]
  assign io_inp_rd_idx_bits = tensorGemm_io_inp_rd_idx_bits; // @[Compute.scala 136:21:@22927.4]
  assign io_wgt_rd_idx_valid = tensorGemm_io_wgt_rd_idx_valid; // @[Compute.scala 137:21:@23445.4]
  assign io_wgt_rd_idx_bits = tensorGemm_io_wgt_rd_idx_bits; // @[Compute.scala 137:21:@23444.4]
  assign io_out_wr_valid = dec_io_isGemm ? tensorGemm_io_out_wr_valid : tensorAlu_io_out_wr_valid; // @[Compute.scala 157:13:@23549.4]
  assign io_out_wr_bits_idx = dec_io_isGemm ? tensorGemm_io_out_wr_bits_idx : tensorAlu_io_out_wr_bits_idx; // @[Compute.scala 157:13:@23548.4]
  assign io_out_wr_bits_data_0_0 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_0 : tensorAlu_io_out_wr_bits_data_0_0; // @[Compute.scala 157:13:@23532.4]
  assign io_out_wr_bits_data_0_1 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_1 : tensorAlu_io_out_wr_bits_data_0_1; // @[Compute.scala 157:13:@23533.4]
  assign io_out_wr_bits_data_0_2 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_2 : tensorAlu_io_out_wr_bits_data_0_2; // @[Compute.scala 157:13:@23534.4]
  assign io_out_wr_bits_data_0_3 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_3 : tensorAlu_io_out_wr_bits_data_0_3; // @[Compute.scala 157:13:@23535.4]
  assign io_out_wr_bits_data_0_4 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_4 : tensorAlu_io_out_wr_bits_data_0_4; // @[Compute.scala 157:13:@23536.4]
  assign io_out_wr_bits_data_0_5 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_5 : tensorAlu_io_out_wr_bits_data_0_5; // @[Compute.scala 157:13:@23537.4]
  assign io_out_wr_bits_data_0_6 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_6 : tensorAlu_io_out_wr_bits_data_0_6; // @[Compute.scala 157:13:@23538.4]
  assign io_out_wr_bits_data_0_7 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_7 : tensorAlu_io_out_wr_bits_data_0_7; // @[Compute.scala 157:13:@23539.4]
  assign io_out_wr_bits_data_0_8 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_8 : tensorAlu_io_out_wr_bits_data_0_8; // @[Compute.scala 157:13:@23540.4]
  assign io_out_wr_bits_data_0_9 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_9 : tensorAlu_io_out_wr_bits_data_0_9; // @[Compute.scala 157:13:@23541.4]
  assign io_out_wr_bits_data_0_10 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_10 : tensorAlu_io_out_wr_bits_data_0_10; // @[Compute.scala 157:13:@23542.4]
  assign io_out_wr_bits_data_0_11 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_11 : tensorAlu_io_out_wr_bits_data_0_11; // @[Compute.scala 157:13:@23543.4]
  assign io_out_wr_bits_data_0_12 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_12 : tensorAlu_io_out_wr_bits_data_0_12; // @[Compute.scala 157:13:@23544.4]
  assign io_out_wr_bits_data_0_13 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_13 : tensorAlu_io_out_wr_bits_data_0_13; // @[Compute.scala 157:13:@23545.4]
  assign io_out_wr_bits_data_0_14 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_14 : tensorAlu_io_out_wr_bits_data_0_14; // @[Compute.scala 157:13:@23546.4]
  assign io_out_wr_bits_data_0_15 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_15 : tensorAlu_io_out_wr_bits_data_0_15; // @[Compute.scala 157:13:@23547.4]
  assign io_finish = _T_7079 & dec_io_isFinish; // @[Compute.scala 168:13:@23575.4]
  assign io_acc_wr_event = tensorAcc_io_tensor_wr_valid; // @[Compute.scala 129:19:@22881.4]
  assign s_0_clock = clock; // @[:@22754.4]
  assign s_0_reset = reset; // @[:@22755.4]
  assign s_0_io_spost = io_i_post_0; // @[Compute.scala 160:17:@23550.4]
  assign s_0_io_swait = dec_io_pop_prev & _T_7083; // @[Compute.scala 162:17:@23555.4]
  assign s_1_clock = clock; // @[:@22757.4]
  assign s_1_reset = reset; // @[:@22758.4]
  assign s_1_io_spost = io_i_post_1; // @[Compute.scala 161:17:@23551.4]
  assign s_1_io_swait = dec_io_pop_next & _T_7083; // @[Compute.scala 163:17:@23559.4]
  assign loadUop_clock = clock; // @[:@22760.4]
  assign loadUop_reset = reset; // @[:@22761.4]
  assign loadUop_io_start = _T_7083 & dec_io_isLoadUop; // @[Compute.scala 116:20:@22833.4]
  assign loadUop_io_inst = inst_q_io_deq_bits; // @[Compute.scala 117:19:@22834.4]
  assign loadUop_io_baddr = io_uop_baddr; // @[Compute.scala 118:20:@22835.4]
  assign loadUop_io_vme_rd_cmd_ready = io_vme_rd_0_cmd_ready; // @[Compute.scala 119:16:@22842.4]
  assign loadUop_io_vme_rd_data_valid = io_vme_rd_0_data_valid; // @[Compute.scala 119:16:@22837.4]
  assign loadUop_io_vme_rd_data_bits = io_vme_rd_0_data_bits; // @[Compute.scala 119:16:@22836.4]
  assign loadUop_io_uop_idx_valid = dec_io_isGemm ? tensorGemm_io_uop_idx_valid : tensorAlu_io_uop_idx_valid; // @[Compute.scala 120:22:@22845.4]
  assign loadUop_io_uop_idx_bits = dec_io_isGemm ? tensorGemm_io_uop_idx_bits : tensorAlu_io_uop_idx_bits; // @[Compute.scala 120:22:@22844.4]
  assign tensorAcc_clock = clock; // @[:@22763.4]
  assign tensorAcc_reset = reset; // @[:@22764.4]
  assign tensorAcc_io_start = _T_7083 & dec_io_isLoadAcc; // @[Compute.scala 123:22:@22849.4]
  assign tensorAcc_io_inst = inst_q_io_deq_bits; // @[Compute.scala 124:21:@22850.4]
  assign tensorAcc_io_baddr = io_acc_baddr; // @[Compute.scala 125:22:@22851.4]
  assign tensorAcc_io_vme_rd_cmd_ready = io_vme_rd_1_cmd_ready; // @[Compute.scala 128:16:@22880.4]
  assign tensorAcc_io_vme_rd_data_valid = io_vme_rd_1_data_valid; // @[Compute.scala 128:16:@22875.4]
  assign tensorAcc_io_vme_rd_data_bits = io_vme_rd_1_data_bits; // @[Compute.scala 128:16:@22874.4]
  assign tensorAcc_io_tensor_rd_idx_valid = dec_io_isGemm ? tensorGemm_io_acc_rd_idx_valid : tensorAlu_io_acc_rd_idx_valid; // @[Compute.scala 126:30:@22854.4]
  assign tensorAcc_io_tensor_rd_idx_bits = dec_io_isGemm ? tensorGemm_io_acc_rd_idx_bits : tensorAlu_io_acc_rd_idx_bits; // @[Compute.scala 126:30:@22853.4]
  assign tensorAcc_io_tensor_wr_valid = dec_io_isGemm ? tensorGemm_io_acc_wr_valid : tensorAlu_io_acc_wr_valid; // @[Compute.scala 127:26:@22873.4]
  assign tensorAcc_io_tensor_wr_bits_idx = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_idx : tensorAlu_io_acc_wr_bits_idx; // @[Compute.scala 127:26:@22872.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_0 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_0 : tensorAlu_io_acc_wr_bits_data_0_0; // @[Compute.scala 127:26:@22856.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_1 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_1 : tensorAlu_io_acc_wr_bits_data_0_1; // @[Compute.scala 127:26:@22857.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_2 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_2 : tensorAlu_io_acc_wr_bits_data_0_2; // @[Compute.scala 127:26:@22858.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_3 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_3 : tensorAlu_io_acc_wr_bits_data_0_3; // @[Compute.scala 127:26:@22859.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_4 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_4 : tensorAlu_io_acc_wr_bits_data_0_4; // @[Compute.scala 127:26:@22860.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_5 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_5 : tensorAlu_io_acc_wr_bits_data_0_5; // @[Compute.scala 127:26:@22861.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_6 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_6 : tensorAlu_io_acc_wr_bits_data_0_6; // @[Compute.scala 127:26:@22862.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_7 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_7 : tensorAlu_io_acc_wr_bits_data_0_7; // @[Compute.scala 127:26:@22863.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_8 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_8 : tensorAlu_io_acc_wr_bits_data_0_8; // @[Compute.scala 127:26:@22864.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_9 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_9 : tensorAlu_io_acc_wr_bits_data_0_9; // @[Compute.scala 127:26:@22865.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_10 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_10 : tensorAlu_io_acc_wr_bits_data_0_10; // @[Compute.scala 127:26:@22866.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_11 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_11 : tensorAlu_io_acc_wr_bits_data_0_11; // @[Compute.scala 127:26:@22867.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_12 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_12 : tensorAlu_io_acc_wr_bits_data_0_12; // @[Compute.scala 127:26:@22868.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_13 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_13 : tensorAlu_io_acc_wr_bits_data_0_13; // @[Compute.scala 127:26:@22869.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_14 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_14 : tensorAlu_io_acc_wr_bits_data_0_14; // @[Compute.scala 127:26:@22870.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_15 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_15 : tensorAlu_io_acc_wr_bits_data_0_15; // @[Compute.scala 127:26:@22871.4]
  assign tensorGemm_clock = clock; // @[:@22766.4]
  assign tensorGemm_reset = reset; // @[:@22767.4]
  assign tensorGemm_io_start = _T_7083 & dec_io_isGemm; // @[Compute.scala 132:23:@22885.4]
  assign tensorGemm_io_inst = inst_q_io_deq_bits; // @[Compute.scala 133:22:@22886.4]
  assign tensorGemm_io_uop_data_valid = loadUop_io_uop_data_valid & dec_io_isGemm; // @[Compute.scala 134:32:@22888.4]
  assign tensorGemm_io_uop_data_bits_u2 = loadUop_io_uop_data_bits_u2; // @[Compute.scala 135:31:@22891.4]
  assign tensorGemm_io_uop_data_bits_u1 = loadUop_io_uop_data_bits_u1; // @[Compute.scala 135:31:@22890.4]
  assign tensorGemm_io_uop_data_bits_u0 = loadUop_io_uop_data_bits_u0; // @[Compute.scala 135:31:@22889.4]
  assign tensorGemm_io_inp_rd_data_valid = io_inp_rd_data_valid; // @[Compute.scala 136:21:@22926.4]
  assign tensorGemm_io_inp_rd_data_bits_0_0 = io_inp_rd_data_bits_0_0; // @[Compute.scala 136:21:@22910.4]
  assign tensorGemm_io_inp_rd_data_bits_0_1 = io_inp_rd_data_bits_0_1; // @[Compute.scala 136:21:@22911.4]
  assign tensorGemm_io_inp_rd_data_bits_0_2 = io_inp_rd_data_bits_0_2; // @[Compute.scala 136:21:@22912.4]
  assign tensorGemm_io_inp_rd_data_bits_0_3 = io_inp_rd_data_bits_0_3; // @[Compute.scala 136:21:@22913.4]
  assign tensorGemm_io_inp_rd_data_bits_0_4 = io_inp_rd_data_bits_0_4; // @[Compute.scala 136:21:@22914.4]
  assign tensorGemm_io_inp_rd_data_bits_0_5 = io_inp_rd_data_bits_0_5; // @[Compute.scala 136:21:@22915.4]
  assign tensorGemm_io_inp_rd_data_bits_0_6 = io_inp_rd_data_bits_0_6; // @[Compute.scala 136:21:@22916.4]
  assign tensorGemm_io_inp_rd_data_bits_0_7 = io_inp_rd_data_bits_0_7; // @[Compute.scala 136:21:@22917.4]
  assign tensorGemm_io_inp_rd_data_bits_0_8 = io_inp_rd_data_bits_0_8; // @[Compute.scala 136:21:@22918.4]
  assign tensorGemm_io_inp_rd_data_bits_0_9 = io_inp_rd_data_bits_0_9; // @[Compute.scala 136:21:@22919.4]
  assign tensorGemm_io_inp_rd_data_bits_0_10 = io_inp_rd_data_bits_0_10; // @[Compute.scala 136:21:@22920.4]
  assign tensorGemm_io_inp_rd_data_bits_0_11 = io_inp_rd_data_bits_0_11; // @[Compute.scala 136:21:@22921.4]
  assign tensorGemm_io_inp_rd_data_bits_0_12 = io_inp_rd_data_bits_0_12; // @[Compute.scala 136:21:@22922.4]
  assign tensorGemm_io_inp_rd_data_bits_0_13 = io_inp_rd_data_bits_0_13; // @[Compute.scala 136:21:@22923.4]
  assign tensorGemm_io_inp_rd_data_bits_0_14 = io_inp_rd_data_bits_0_14; // @[Compute.scala 136:21:@22924.4]
  assign tensorGemm_io_inp_rd_data_bits_0_15 = io_inp_rd_data_bits_0_15; // @[Compute.scala 136:21:@22925.4]
  assign tensorGemm_io_wgt_rd_data_valid = io_wgt_rd_data_valid; // @[Compute.scala 137:21:@23443.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_0 = io_wgt_rd_data_bits_0_0; // @[Compute.scala 137:21:@23187.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_1 = io_wgt_rd_data_bits_0_1; // @[Compute.scala 137:21:@23188.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_2 = io_wgt_rd_data_bits_0_2; // @[Compute.scala 137:21:@23189.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_3 = io_wgt_rd_data_bits_0_3; // @[Compute.scala 137:21:@23190.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_4 = io_wgt_rd_data_bits_0_4; // @[Compute.scala 137:21:@23191.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_5 = io_wgt_rd_data_bits_0_5; // @[Compute.scala 137:21:@23192.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_6 = io_wgt_rd_data_bits_0_6; // @[Compute.scala 137:21:@23193.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_7 = io_wgt_rd_data_bits_0_7; // @[Compute.scala 137:21:@23194.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_8 = io_wgt_rd_data_bits_0_8; // @[Compute.scala 137:21:@23195.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_9 = io_wgt_rd_data_bits_0_9; // @[Compute.scala 137:21:@23196.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_10 = io_wgt_rd_data_bits_0_10; // @[Compute.scala 137:21:@23197.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_11 = io_wgt_rd_data_bits_0_11; // @[Compute.scala 137:21:@23198.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_12 = io_wgt_rd_data_bits_0_12; // @[Compute.scala 137:21:@23199.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_13 = io_wgt_rd_data_bits_0_13; // @[Compute.scala 137:21:@23200.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_14 = io_wgt_rd_data_bits_0_14; // @[Compute.scala 137:21:@23201.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_15 = io_wgt_rd_data_bits_0_15; // @[Compute.scala 137:21:@23202.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_0 = io_wgt_rd_data_bits_1_0; // @[Compute.scala 137:21:@23203.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_1 = io_wgt_rd_data_bits_1_1; // @[Compute.scala 137:21:@23204.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_2 = io_wgt_rd_data_bits_1_2; // @[Compute.scala 137:21:@23205.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_3 = io_wgt_rd_data_bits_1_3; // @[Compute.scala 137:21:@23206.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_4 = io_wgt_rd_data_bits_1_4; // @[Compute.scala 137:21:@23207.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_5 = io_wgt_rd_data_bits_1_5; // @[Compute.scala 137:21:@23208.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_6 = io_wgt_rd_data_bits_1_6; // @[Compute.scala 137:21:@23209.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_7 = io_wgt_rd_data_bits_1_7; // @[Compute.scala 137:21:@23210.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_8 = io_wgt_rd_data_bits_1_8; // @[Compute.scala 137:21:@23211.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_9 = io_wgt_rd_data_bits_1_9; // @[Compute.scala 137:21:@23212.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_10 = io_wgt_rd_data_bits_1_10; // @[Compute.scala 137:21:@23213.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_11 = io_wgt_rd_data_bits_1_11; // @[Compute.scala 137:21:@23214.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_12 = io_wgt_rd_data_bits_1_12; // @[Compute.scala 137:21:@23215.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_13 = io_wgt_rd_data_bits_1_13; // @[Compute.scala 137:21:@23216.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_14 = io_wgt_rd_data_bits_1_14; // @[Compute.scala 137:21:@23217.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_15 = io_wgt_rd_data_bits_1_15; // @[Compute.scala 137:21:@23218.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_0 = io_wgt_rd_data_bits_2_0; // @[Compute.scala 137:21:@23219.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_1 = io_wgt_rd_data_bits_2_1; // @[Compute.scala 137:21:@23220.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_2 = io_wgt_rd_data_bits_2_2; // @[Compute.scala 137:21:@23221.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_3 = io_wgt_rd_data_bits_2_3; // @[Compute.scala 137:21:@23222.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_4 = io_wgt_rd_data_bits_2_4; // @[Compute.scala 137:21:@23223.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_5 = io_wgt_rd_data_bits_2_5; // @[Compute.scala 137:21:@23224.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_6 = io_wgt_rd_data_bits_2_6; // @[Compute.scala 137:21:@23225.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_7 = io_wgt_rd_data_bits_2_7; // @[Compute.scala 137:21:@23226.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_8 = io_wgt_rd_data_bits_2_8; // @[Compute.scala 137:21:@23227.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_9 = io_wgt_rd_data_bits_2_9; // @[Compute.scala 137:21:@23228.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_10 = io_wgt_rd_data_bits_2_10; // @[Compute.scala 137:21:@23229.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_11 = io_wgt_rd_data_bits_2_11; // @[Compute.scala 137:21:@23230.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_12 = io_wgt_rd_data_bits_2_12; // @[Compute.scala 137:21:@23231.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_13 = io_wgt_rd_data_bits_2_13; // @[Compute.scala 137:21:@23232.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_14 = io_wgt_rd_data_bits_2_14; // @[Compute.scala 137:21:@23233.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_15 = io_wgt_rd_data_bits_2_15; // @[Compute.scala 137:21:@23234.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_0 = io_wgt_rd_data_bits_3_0; // @[Compute.scala 137:21:@23235.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_1 = io_wgt_rd_data_bits_3_1; // @[Compute.scala 137:21:@23236.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_2 = io_wgt_rd_data_bits_3_2; // @[Compute.scala 137:21:@23237.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_3 = io_wgt_rd_data_bits_3_3; // @[Compute.scala 137:21:@23238.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_4 = io_wgt_rd_data_bits_3_4; // @[Compute.scala 137:21:@23239.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_5 = io_wgt_rd_data_bits_3_5; // @[Compute.scala 137:21:@23240.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_6 = io_wgt_rd_data_bits_3_6; // @[Compute.scala 137:21:@23241.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_7 = io_wgt_rd_data_bits_3_7; // @[Compute.scala 137:21:@23242.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_8 = io_wgt_rd_data_bits_3_8; // @[Compute.scala 137:21:@23243.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_9 = io_wgt_rd_data_bits_3_9; // @[Compute.scala 137:21:@23244.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_10 = io_wgt_rd_data_bits_3_10; // @[Compute.scala 137:21:@23245.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_11 = io_wgt_rd_data_bits_3_11; // @[Compute.scala 137:21:@23246.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_12 = io_wgt_rd_data_bits_3_12; // @[Compute.scala 137:21:@23247.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_13 = io_wgt_rd_data_bits_3_13; // @[Compute.scala 137:21:@23248.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_14 = io_wgt_rd_data_bits_3_14; // @[Compute.scala 137:21:@23249.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_15 = io_wgt_rd_data_bits_3_15; // @[Compute.scala 137:21:@23250.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_0 = io_wgt_rd_data_bits_4_0; // @[Compute.scala 137:21:@23251.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_1 = io_wgt_rd_data_bits_4_1; // @[Compute.scala 137:21:@23252.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_2 = io_wgt_rd_data_bits_4_2; // @[Compute.scala 137:21:@23253.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_3 = io_wgt_rd_data_bits_4_3; // @[Compute.scala 137:21:@23254.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_4 = io_wgt_rd_data_bits_4_4; // @[Compute.scala 137:21:@23255.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_5 = io_wgt_rd_data_bits_4_5; // @[Compute.scala 137:21:@23256.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_6 = io_wgt_rd_data_bits_4_6; // @[Compute.scala 137:21:@23257.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_7 = io_wgt_rd_data_bits_4_7; // @[Compute.scala 137:21:@23258.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_8 = io_wgt_rd_data_bits_4_8; // @[Compute.scala 137:21:@23259.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_9 = io_wgt_rd_data_bits_4_9; // @[Compute.scala 137:21:@23260.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_10 = io_wgt_rd_data_bits_4_10; // @[Compute.scala 137:21:@23261.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_11 = io_wgt_rd_data_bits_4_11; // @[Compute.scala 137:21:@23262.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_12 = io_wgt_rd_data_bits_4_12; // @[Compute.scala 137:21:@23263.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_13 = io_wgt_rd_data_bits_4_13; // @[Compute.scala 137:21:@23264.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_14 = io_wgt_rd_data_bits_4_14; // @[Compute.scala 137:21:@23265.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_15 = io_wgt_rd_data_bits_4_15; // @[Compute.scala 137:21:@23266.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_0 = io_wgt_rd_data_bits_5_0; // @[Compute.scala 137:21:@23267.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_1 = io_wgt_rd_data_bits_5_1; // @[Compute.scala 137:21:@23268.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_2 = io_wgt_rd_data_bits_5_2; // @[Compute.scala 137:21:@23269.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_3 = io_wgt_rd_data_bits_5_3; // @[Compute.scala 137:21:@23270.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_4 = io_wgt_rd_data_bits_5_4; // @[Compute.scala 137:21:@23271.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_5 = io_wgt_rd_data_bits_5_5; // @[Compute.scala 137:21:@23272.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_6 = io_wgt_rd_data_bits_5_6; // @[Compute.scala 137:21:@23273.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_7 = io_wgt_rd_data_bits_5_7; // @[Compute.scala 137:21:@23274.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_8 = io_wgt_rd_data_bits_5_8; // @[Compute.scala 137:21:@23275.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_9 = io_wgt_rd_data_bits_5_9; // @[Compute.scala 137:21:@23276.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_10 = io_wgt_rd_data_bits_5_10; // @[Compute.scala 137:21:@23277.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_11 = io_wgt_rd_data_bits_5_11; // @[Compute.scala 137:21:@23278.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_12 = io_wgt_rd_data_bits_5_12; // @[Compute.scala 137:21:@23279.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_13 = io_wgt_rd_data_bits_5_13; // @[Compute.scala 137:21:@23280.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_14 = io_wgt_rd_data_bits_5_14; // @[Compute.scala 137:21:@23281.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_15 = io_wgt_rd_data_bits_5_15; // @[Compute.scala 137:21:@23282.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_0 = io_wgt_rd_data_bits_6_0; // @[Compute.scala 137:21:@23283.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_1 = io_wgt_rd_data_bits_6_1; // @[Compute.scala 137:21:@23284.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_2 = io_wgt_rd_data_bits_6_2; // @[Compute.scala 137:21:@23285.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_3 = io_wgt_rd_data_bits_6_3; // @[Compute.scala 137:21:@23286.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_4 = io_wgt_rd_data_bits_6_4; // @[Compute.scala 137:21:@23287.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_5 = io_wgt_rd_data_bits_6_5; // @[Compute.scala 137:21:@23288.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_6 = io_wgt_rd_data_bits_6_6; // @[Compute.scala 137:21:@23289.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_7 = io_wgt_rd_data_bits_6_7; // @[Compute.scala 137:21:@23290.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_8 = io_wgt_rd_data_bits_6_8; // @[Compute.scala 137:21:@23291.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_9 = io_wgt_rd_data_bits_6_9; // @[Compute.scala 137:21:@23292.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_10 = io_wgt_rd_data_bits_6_10; // @[Compute.scala 137:21:@23293.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_11 = io_wgt_rd_data_bits_6_11; // @[Compute.scala 137:21:@23294.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_12 = io_wgt_rd_data_bits_6_12; // @[Compute.scala 137:21:@23295.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_13 = io_wgt_rd_data_bits_6_13; // @[Compute.scala 137:21:@23296.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_14 = io_wgt_rd_data_bits_6_14; // @[Compute.scala 137:21:@23297.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_15 = io_wgt_rd_data_bits_6_15; // @[Compute.scala 137:21:@23298.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_0 = io_wgt_rd_data_bits_7_0; // @[Compute.scala 137:21:@23299.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_1 = io_wgt_rd_data_bits_7_1; // @[Compute.scala 137:21:@23300.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_2 = io_wgt_rd_data_bits_7_2; // @[Compute.scala 137:21:@23301.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_3 = io_wgt_rd_data_bits_7_3; // @[Compute.scala 137:21:@23302.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_4 = io_wgt_rd_data_bits_7_4; // @[Compute.scala 137:21:@23303.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_5 = io_wgt_rd_data_bits_7_5; // @[Compute.scala 137:21:@23304.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_6 = io_wgt_rd_data_bits_7_6; // @[Compute.scala 137:21:@23305.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_7 = io_wgt_rd_data_bits_7_7; // @[Compute.scala 137:21:@23306.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_8 = io_wgt_rd_data_bits_7_8; // @[Compute.scala 137:21:@23307.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_9 = io_wgt_rd_data_bits_7_9; // @[Compute.scala 137:21:@23308.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_10 = io_wgt_rd_data_bits_7_10; // @[Compute.scala 137:21:@23309.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_11 = io_wgt_rd_data_bits_7_11; // @[Compute.scala 137:21:@23310.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_12 = io_wgt_rd_data_bits_7_12; // @[Compute.scala 137:21:@23311.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_13 = io_wgt_rd_data_bits_7_13; // @[Compute.scala 137:21:@23312.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_14 = io_wgt_rd_data_bits_7_14; // @[Compute.scala 137:21:@23313.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_15 = io_wgt_rd_data_bits_7_15; // @[Compute.scala 137:21:@23314.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_0 = io_wgt_rd_data_bits_8_0; // @[Compute.scala 137:21:@23315.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_1 = io_wgt_rd_data_bits_8_1; // @[Compute.scala 137:21:@23316.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_2 = io_wgt_rd_data_bits_8_2; // @[Compute.scala 137:21:@23317.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_3 = io_wgt_rd_data_bits_8_3; // @[Compute.scala 137:21:@23318.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_4 = io_wgt_rd_data_bits_8_4; // @[Compute.scala 137:21:@23319.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_5 = io_wgt_rd_data_bits_8_5; // @[Compute.scala 137:21:@23320.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_6 = io_wgt_rd_data_bits_8_6; // @[Compute.scala 137:21:@23321.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_7 = io_wgt_rd_data_bits_8_7; // @[Compute.scala 137:21:@23322.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_8 = io_wgt_rd_data_bits_8_8; // @[Compute.scala 137:21:@23323.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_9 = io_wgt_rd_data_bits_8_9; // @[Compute.scala 137:21:@23324.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_10 = io_wgt_rd_data_bits_8_10; // @[Compute.scala 137:21:@23325.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_11 = io_wgt_rd_data_bits_8_11; // @[Compute.scala 137:21:@23326.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_12 = io_wgt_rd_data_bits_8_12; // @[Compute.scala 137:21:@23327.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_13 = io_wgt_rd_data_bits_8_13; // @[Compute.scala 137:21:@23328.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_14 = io_wgt_rd_data_bits_8_14; // @[Compute.scala 137:21:@23329.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_15 = io_wgt_rd_data_bits_8_15; // @[Compute.scala 137:21:@23330.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_0 = io_wgt_rd_data_bits_9_0; // @[Compute.scala 137:21:@23331.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_1 = io_wgt_rd_data_bits_9_1; // @[Compute.scala 137:21:@23332.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_2 = io_wgt_rd_data_bits_9_2; // @[Compute.scala 137:21:@23333.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_3 = io_wgt_rd_data_bits_9_3; // @[Compute.scala 137:21:@23334.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_4 = io_wgt_rd_data_bits_9_4; // @[Compute.scala 137:21:@23335.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_5 = io_wgt_rd_data_bits_9_5; // @[Compute.scala 137:21:@23336.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_6 = io_wgt_rd_data_bits_9_6; // @[Compute.scala 137:21:@23337.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_7 = io_wgt_rd_data_bits_9_7; // @[Compute.scala 137:21:@23338.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_8 = io_wgt_rd_data_bits_9_8; // @[Compute.scala 137:21:@23339.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_9 = io_wgt_rd_data_bits_9_9; // @[Compute.scala 137:21:@23340.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_10 = io_wgt_rd_data_bits_9_10; // @[Compute.scala 137:21:@23341.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_11 = io_wgt_rd_data_bits_9_11; // @[Compute.scala 137:21:@23342.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_12 = io_wgt_rd_data_bits_9_12; // @[Compute.scala 137:21:@23343.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_13 = io_wgt_rd_data_bits_9_13; // @[Compute.scala 137:21:@23344.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_14 = io_wgt_rd_data_bits_9_14; // @[Compute.scala 137:21:@23345.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_15 = io_wgt_rd_data_bits_9_15; // @[Compute.scala 137:21:@23346.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_0 = io_wgt_rd_data_bits_10_0; // @[Compute.scala 137:21:@23347.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_1 = io_wgt_rd_data_bits_10_1; // @[Compute.scala 137:21:@23348.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_2 = io_wgt_rd_data_bits_10_2; // @[Compute.scala 137:21:@23349.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_3 = io_wgt_rd_data_bits_10_3; // @[Compute.scala 137:21:@23350.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_4 = io_wgt_rd_data_bits_10_4; // @[Compute.scala 137:21:@23351.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_5 = io_wgt_rd_data_bits_10_5; // @[Compute.scala 137:21:@23352.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_6 = io_wgt_rd_data_bits_10_6; // @[Compute.scala 137:21:@23353.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_7 = io_wgt_rd_data_bits_10_7; // @[Compute.scala 137:21:@23354.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_8 = io_wgt_rd_data_bits_10_8; // @[Compute.scala 137:21:@23355.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_9 = io_wgt_rd_data_bits_10_9; // @[Compute.scala 137:21:@23356.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_10 = io_wgt_rd_data_bits_10_10; // @[Compute.scala 137:21:@23357.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_11 = io_wgt_rd_data_bits_10_11; // @[Compute.scala 137:21:@23358.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_12 = io_wgt_rd_data_bits_10_12; // @[Compute.scala 137:21:@23359.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_13 = io_wgt_rd_data_bits_10_13; // @[Compute.scala 137:21:@23360.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_14 = io_wgt_rd_data_bits_10_14; // @[Compute.scala 137:21:@23361.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_15 = io_wgt_rd_data_bits_10_15; // @[Compute.scala 137:21:@23362.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_0 = io_wgt_rd_data_bits_11_0; // @[Compute.scala 137:21:@23363.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_1 = io_wgt_rd_data_bits_11_1; // @[Compute.scala 137:21:@23364.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_2 = io_wgt_rd_data_bits_11_2; // @[Compute.scala 137:21:@23365.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_3 = io_wgt_rd_data_bits_11_3; // @[Compute.scala 137:21:@23366.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_4 = io_wgt_rd_data_bits_11_4; // @[Compute.scala 137:21:@23367.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_5 = io_wgt_rd_data_bits_11_5; // @[Compute.scala 137:21:@23368.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_6 = io_wgt_rd_data_bits_11_6; // @[Compute.scala 137:21:@23369.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_7 = io_wgt_rd_data_bits_11_7; // @[Compute.scala 137:21:@23370.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_8 = io_wgt_rd_data_bits_11_8; // @[Compute.scala 137:21:@23371.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_9 = io_wgt_rd_data_bits_11_9; // @[Compute.scala 137:21:@23372.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_10 = io_wgt_rd_data_bits_11_10; // @[Compute.scala 137:21:@23373.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_11 = io_wgt_rd_data_bits_11_11; // @[Compute.scala 137:21:@23374.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_12 = io_wgt_rd_data_bits_11_12; // @[Compute.scala 137:21:@23375.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_13 = io_wgt_rd_data_bits_11_13; // @[Compute.scala 137:21:@23376.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_14 = io_wgt_rd_data_bits_11_14; // @[Compute.scala 137:21:@23377.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_15 = io_wgt_rd_data_bits_11_15; // @[Compute.scala 137:21:@23378.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_0 = io_wgt_rd_data_bits_12_0; // @[Compute.scala 137:21:@23379.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_1 = io_wgt_rd_data_bits_12_1; // @[Compute.scala 137:21:@23380.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_2 = io_wgt_rd_data_bits_12_2; // @[Compute.scala 137:21:@23381.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_3 = io_wgt_rd_data_bits_12_3; // @[Compute.scala 137:21:@23382.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_4 = io_wgt_rd_data_bits_12_4; // @[Compute.scala 137:21:@23383.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_5 = io_wgt_rd_data_bits_12_5; // @[Compute.scala 137:21:@23384.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_6 = io_wgt_rd_data_bits_12_6; // @[Compute.scala 137:21:@23385.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_7 = io_wgt_rd_data_bits_12_7; // @[Compute.scala 137:21:@23386.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_8 = io_wgt_rd_data_bits_12_8; // @[Compute.scala 137:21:@23387.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_9 = io_wgt_rd_data_bits_12_9; // @[Compute.scala 137:21:@23388.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_10 = io_wgt_rd_data_bits_12_10; // @[Compute.scala 137:21:@23389.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_11 = io_wgt_rd_data_bits_12_11; // @[Compute.scala 137:21:@23390.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_12 = io_wgt_rd_data_bits_12_12; // @[Compute.scala 137:21:@23391.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_13 = io_wgt_rd_data_bits_12_13; // @[Compute.scala 137:21:@23392.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_14 = io_wgt_rd_data_bits_12_14; // @[Compute.scala 137:21:@23393.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_15 = io_wgt_rd_data_bits_12_15; // @[Compute.scala 137:21:@23394.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_0 = io_wgt_rd_data_bits_13_0; // @[Compute.scala 137:21:@23395.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_1 = io_wgt_rd_data_bits_13_1; // @[Compute.scala 137:21:@23396.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_2 = io_wgt_rd_data_bits_13_2; // @[Compute.scala 137:21:@23397.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_3 = io_wgt_rd_data_bits_13_3; // @[Compute.scala 137:21:@23398.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_4 = io_wgt_rd_data_bits_13_4; // @[Compute.scala 137:21:@23399.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_5 = io_wgt_rd_data_bits_13_5; // @[Compute.scala 137:21:@23400.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_6 = io_wgt_rd_data_bits_13_6; // @[Compute.scala 137:21:@23401.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_7 = io_wgt_rd_data_bits_13_7; // @[Compute.scala 137:21:@23402.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_8 = io_wgt_rd_data_bits_13_8; // @[Compute.scala 137:21:@23403.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_9 = io_wgt_rd_data_bits_13_9; // @[Compute.scala 137:21:@23404.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_10 = io_wgt_rd_data_bits_13_10; // @[Compute.scala 137:21:@23405.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_11 = io_wgt_rd_data_bits_13_11; // @[Compute.scala 137:21:@23406.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_12 = io_wgt_rd_data_bits_13_12; // @[Compute.scala 137:21:@23407.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_13 = io_wgt_rd_data_bits_13_13; // @[Compute.scala 137:21:@23408.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_14 = io_wgt_rd_data_bits_13_14; // @[Compute.scala 137:21:@23409.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_15 = io_wgt_rd_data_bits_13_15; // @[Compute.scala 137:21:@23410.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_0 = io_wgt_rd_data_bits_14_0; // @[Compute.scala 137:21:@23411.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_1 = io_wgt_rd_data_bits_14_1; // @[Compute.scala 137:21:@23412.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_2 = io_wgt_rd_data_bits_14_2; // @[Compute.scala 137:21:@23413.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_3 = io_wgt_rd_data_bits_14_3; // @[Compute.scala 137:21:@23414.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_4 = io_wgt_rd_data_bits_14_4; // @[Compute.scala 137:21:@23415.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_5 = io_wgt_rd_data_bits_14_5; // @[Compute.scala 137:21:@23416.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_6 = io_wgt_rd_data_bits_14_6; // @[Compute.scala 137:21:@23417.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_7 = io_wgt_rd_data_bits_14_7; // @[Compute.scala 137:21:@23418.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_8 = io_wgt_rd_data_bits_14_8; // @[Compute.scala 137:21:@23419.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_9 = io_wgt_rd_data_bits_14_9; // @[Compute.scala 137:21:@23420.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_10 = io_wgt_rd_data_bits_14_10; // @[Compute.scala 137:21:@23421.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_11 = io_wgt_rd_data_bits_14_11; // @[Compute.scala 137:21:@23422.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_12 = io_wgt_rd_data_bits_14_12; // @[Compute.scala 137:21:@23423.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_13 = io_wgt_rd_data_bits_14_13; // @[Compute.scala 137:21:@23424.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_14 = io_wgt_rd_data_bits_14_14; // @[Compute.scala 137:21:@23425.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_15 = io_wgt_rd_data_bits_14_15; // @[Compute.scala 137:21:@23426.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_0 = io_wgt_rd_data_bits_15_0; // @[Compute.scala 137:21:@23427.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_1 = io_wgt_rd_data_bits_15_1; // @[Compute.scala 137:21:@23428.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_2 = io_wgt_rd_data_bits_15_2; // @[Compute.scala 137:21:@23429.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_3 = io_wgt_rd_data_bits_15_3; // @[Compute.scala 137:21:@23430.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_4 = io_wgt_rd_data_bits_15_4; // @[Compute.scala 137:21:@23431.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_5 = io_wgt_rd_data_bits_15_5; // @[Compute.scala 137:21:@23432.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_6 = io_wgt_rd_data_bits_15_6; // @[Compute.scala 137:21:@23433.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_7 = io_wgt_rd_data_bits_15_7; // @[Compute.scala 137:21:@23434.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_8 = io_wgt_rd_data_bits_15_8; // @[Compute.scala 137:21:@23435.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_9 = io_wgt_rd_data_bits_15_9; // @[Compute.scala 137:21:@23436.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_10 = io_wgt_rd_data_bits_15_10; // @[Compute.scala 137:21:@23437.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_11 = io_wgt_rd_data_bits_15_11; // @[Compute.scala 137:21:@23438.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_12 = io_wgt_rd_data_bits_15_12; // @[Compute.scala 137:21:@23439.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_13 = io_wgt_rd_data_bits_15_13; // @[Compute.scala 137:21:@23440.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_14 = io_wgt_rd_data_bits_15_14; // @[Compute.scala 137:21:@23441.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_15 = io_wgt_rd_data_bits_15_15; // @[Compute.scala 137:21:@23442.4]
  assign tensorGemm_io_acc_rd_data_valid = tensorAcc_io_tensor_rd_data_valid & dec_io_isGemm; // @[Compute.scala 138:35:@23447.4]
  assign tensorGemm_io_acc_rd_data_bits_0_0 = tensorAcc_io_tensor_rd_data_bits_0_0; // @[Compute.scala 139:34:@23448.4]
  assign tensorGemm_io_acc_rd_data_bits_0_1 = tensorAcc_io_tensor_rd_data_bits_0_1; // @[Compute.scala 139:34:@23449.4]
  assign tensorGemm_io_acc_rd_data_bits_0_2 = tensorAcc_io_tensor_rd_data_bits_0_2; // @[Compute.scala 139:34:@23450.4]
  assign tensorGemm_io_acc_rd_data_bits_0_3 = tensorAcc_io_tensor_rd_data_bits_0_3; // @[Compute.scala 139:34:@23451.4]
  assign tensorGemm_io_acc_rd_data_bits_0_4 = tensorAcc_io_tensor_rd_data_bits_0_4; // @[Compute.scala 139:34:@23452.4]
  assign tensorGemm_io_acc_rd_data_bits_0_5 = tensorAcc_io_tensor_rd_data_bits_0_5; // @[Compute.scala 139:34:@23453.4]
  assign tensorGemm_io_acc_rd_data_bits_0_6 = tensorAcc_io_tensor_rd_data_bits_0_6; // @[Compute.scala 139:34:@23454.4]
  assign tensorGemm_io_acc_rd_data_bits_0_7 = tensorAcc_io_tensor_rd_data_bits_0_7; // @[Compute.scala 139:34:@23455.4]
  assign tensorGemm_io_acc_rd_data_bits_0_8 = tensorAcc_io_tensor_rd_data_bits_0_8; // @[Compute.scala 139:34:@23456.4]
  assign tensorGemm_io_acc_rd_data_bits_0_9 = tensorAcc_io_tensor_rd_data_bits_0_9; // @[Compute.scala 139:34:@23457.4]
  assign tensorGemm_io_acc_rd_data_bits_0_10 = tensorAcc_io_tensor_rd_data_bits_0_10; // @[Compute.scala 139:34:@23458.4]
  assign tensorGemm_io_acc_rd_data_bits_0_11 = tensorAcc_io_tensor_rd_data_bits_0_11; // @[Compute.scala 139:34:@23459.4]
  assign tensorGemm_io_acc_rd_data_bits_0_12 = tensorAcc_io_tensor_rd_data_bits_0_12; // @[Compute.scala 139:34:@23460.4]
  assign tensorGemm_io_acc_rd_data_bits_0_13 = tensorAcc_io_tensor_rd_data_bits_0_13; // @[Compute.scala 139:34:@23461.4]
  assign tensorGemm_io_acc_rd_data_bits_0_14 = tensorAcc_io_tensor_rd_data_bits_0_14; // @[Compute.scala 139:34:@23462.4]
  assign tensorGemm_io_acc_rd_data_bits_0_15 = tensorAcc_io_tensor_rd_data_bits_0_15; // @[Compute.scala 139:34:@23463.4]
  assign tensorAlu_clock = clock; // @[:@22769.4]
  assign tensorAlu_reset = reset; // @[:@22770.4]
  assign tensorAlu_io_start = _T_7083 & dec_io_isAlu; // @[Compute.scala 144:22:@23485.4]
  assign tensorAlu_io_inst = inst_q_io_deq_bits; // @[Compute.scala 145:21:@23486.4]
  assign tensorAlu_io_uop_data_valid = loadUop_io_uop_data_valid & dec_io_isAlu; // @[Compute.scala 146:31:@23488.4]
  assign tensorAlu_io_uop_data_bits_u1 = loadUop_io_uop_data_bits_u1; // @[Compute.scala 147:30:@23490.4]
  assign tensorAlu_io_uop_data_bits_u0 = loadUop_io_uop_data_bits_u0; // @[Compute.scala 147:30:@23489.4]
  assign tensorAlu_io_acc_rd_data_valid = tensorAcc_io_tensor_rd_data_valid & dec_io_isAlu; // @[Compute.scala 148:34:@23493.4]
  assign tensorAlu_io_acc_rd_data_bits_0_0 = tensorAcc_io_tensor_rd_data_bits_0_0; // @[Compute.scala 149:33:@23494.4]
  assign tensorAlu_io_acc_rd_data_bits_0_1 = tensorAcc_io_tensor_rd_data_bits_0_1; // @[Compute.scala 149:33:@23495.4]
  assign tensorAlu_io_acc_rd_data_bits_0_2 = tensorAcc_io_tensor_rd_data_bits_0_2; // @[Compute.scala 149:33:@23496.4]
  assign tensorAlu_io_acc_rd_data_bits_0_3 = tensorAcc_io_tensor_rd_data_bits_0_3; // @[Compute.scala 149:33:@23497.4]
  assign tensorAlu_io_acc_rd_data_bits_0_4 = tensorAcc_io_tensor_rd_data_bits_0_4; // @[Compute.scala 149:33:@23498.4]
  assign tensorAlu_io_acc_rd_data_bits_0_5 = tensorAcc_io_tensor_rd_data_bits_0_5; // @[Compute.scala 149:33:@23499.4]
  assign tensorAlu_io_acc_rd_data_bits_0_6 = tensorAcc_io_tensor_rd_data_bits_0_6; // @[Compute.scala 149:33:@23500.4]
  assign tensorAlu_io_acc_rd_data_bits_0_7 = tensorAcc_io_tensor_rd_data_bits_0_7; // @[Compute.scala 149:33:@23501.4]
  assign tensorAlu_io_acc_rd_data_bits_0_8 = tensorAcc_io_tensor_rd_data_bits_0_8; // @[Compute.scala 149:33:@23502.4]
  assign tensorAlu_io_acc_rd_data_bits_0_9 = tensorAcc_io_tensor_rd_data_bits_0_9; // @[Compute.scala 149:33:@23503.4]
  assign tensorAlu_io_acc_rd_data_bits_0_10 = tensorAcc_io_tensor_rd_data_bits_0_10; // @[Compute.scala 149:33:@23504.4]
  assign tensorAlu_io_acc_rd_data_bits_0_11 = tensorAcc_io_tensor_rd_data_bits_0_11; // @[Compute.scala 149:33:@23505.4]
  assign tensorAlu_io_acc_rd_data_bits_0_12 = tensorAcc_io_tensor_rd_data_bits_0_12; // @[Compute.scala 149:33:@23506.4]
  assign tensorAlu_io_acc_rd_data_bits_0_13 = tensorAcc_io_tensor_rd_data_bits_0_13; // @[Compute.scala 149:33:@23507.4]
  assign tensorAlu_io_acc_rd_data_bits_0_14 = tensorAcc_io_tensor_rd_data_bits_0_14; // @[Compute.scala 149:33:@23508.4]
  assign tensorAlu_io_acc_rd_data_bits_0_15 = tensorAcc_io_tensor_rd_data_bits_0_15; // @[Compute.scala 149:33:@23509.4]
  assign inst_q_clock = clock; // @[:@22772.4]
  assign inst_q_reset = reset; // @[:@22773.4]
  assign inst_q_io_enq_valid = io_inst_valid; // @[Compute.scala 112:17:@22823.4]
  assign inst_q_io_enq_bits = io_inst_bits; // @[Compute.scala 112:17:@22822.4]
  assign inst_q_io_deq_ready = _T_7079 | _T_7080; // @[Compute.scala 113:23:@22829.4]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Compute.scala 65:15:@22777.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_7073) begin
        if (start) begin
          if (dec_io_isSync) begin
            state <= 2'h1;
          end else begin
            if (_T_7075) begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_7076) begin
          state <= 2'h0;
        end else begin
          if (_T_7077) begin
            if (done) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module StoreDecode( // @[:@23656.2]
  input  [127:0] io_inst, // @[:@23659.4]
  output         io_push_prev, // @[:@23659.4]
  output         io_pop_prev, // @[:@23659.4]
  output         io_isStore, // @[:@23659.4]
  output         io_isSync // @[:@23659.4]
);
  wire [15:0] dec_xsize; // @[Decode.scala 225:29:@23684.4]
  wire [127:0] _T_37; // @[Decode.scala 228:25:@23698.4]
  wire  _T_38; // @[Decode.scala 228:25:@23699.4]
  wire  _T_40; // @[Decode.scala 228:46:@23700.4]
  wire  _T_47; // @[Decode.scala 229:45:@23705.4]
  assign dec_xsize = io_inst[95:80]; // @[Decode.scala 225:29:@23684.4]
  assign _T_37 = io_inst & 128'h7; // @[Decode.scala 228:25:@23698.4]
  assign _T_38 = 128'h1 == _T_37; // @[Decode.scala 228:25:@23699.4]
  assign _T_40 = dec_xsize != 16'h0; // @[Decode.scala 228:46:@23700.4]
  assign _T_47 = dec_xsize == 16'h0; // @[Decode.scala 229:45:@23705.4]
  assign io_push_prev = io_inst[5]; // @[Decode.scala 226:16:@23696.4]
  assign io_pop_prev = io_inst[3]; // @[Decode.scala 227:15:@23697.4]
  assign io_isStore = _T_38 & _T_40; // @[Decode.scala 228:14:@23702.4]
  assign io_isSync = _T_38 & _T_47; // @[Decode.scala 229:13:@23707.4]
endmodule
module TensorStore( // @[:@23709.2]
  input          clock, // @[:@23710.4]
  input          reset, // @[:@23711.4]
  input          io_start, // @[:@23712.4]
  output         io_done, // @[:@23712.4]
  input  [127:0] io_inst, // @[:@23712.4]
  input  [31:0]  io_baddr, // @[:@23712.4]
  input          io_vme_wr_cmd_ready, // @[:@23712.4]
  output         io_vme_wr_cmd_valid, // @[:@23712.4]
  output [31:0]  io_vme_wr_cmd_bits_addr, // @[:@23712.4]
  output [7:0]   io_vme_wr_cmd_bits_len, // @[:@23712.4]
  input          io_vme_wr_data_ready, // @[:@23712.4]
  output         io_vme_wr_data_valid, // @[:@23712.4]
  output [63:0]  io_vme_wr_data_bits, // @[:@23712.4]
  input          io_vme_wr_ack, // @[:@23712.4]
  input          io_tensor_wr_valid, // @[:@23712.4]
  input  [10:0]  io_tensor_wr_bits_idx, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_0, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_1, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_2, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_3, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_4, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_5, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_6, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_7, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_8, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_9, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_10, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_11, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_12, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_13, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_14, // @[:@23712.4]
  input  [7:0]   io_tensor_wr_bits_data_0_15 // @[:@23712.4]
);
  reg [63:0] tensorFile_0_0 [0:2047]; // @[TensorStore.scala 152:16:@23954.4]
  reg [63:0] _RAND_0;
  wire [63:0] tensorFile_0_0__T_914_data; // @[TensorStore.scala 152:16:@23954.4]
  wire [10:0] tensorFile_0_0__T_914_addr; // @[TensorStore.scala 152:16:@23954.4]
  wire [63:0] tensorFile_0_0__T_836_data; // @[TensorStore.scala 152:16:@23954.4]
  wire [10:0] tensorFile_0_0__T_836_addr; // @[TensorStore.scala 152:16:@23954.4]
  wire  tensorFile_0_0__T_836_mask; // @[TensorStore.scala 152:16:@23954.4]
  wire  tensorFile_0_0__T_836_en; // @[TensorStore.scala 152:16:@23954.4]
  reg [63:0] tensorFile_0_1 [0:2047]; // @[TensorStore.scala 152:16:@23954.4]
  reg [63:0] _RAND_1;
  wire [63:0] tensorFile_0_1__T_914_data; // @[TensorStore.scala 152:16:@23954.4]
  wire [10:0] tensorFile_0_1__T_914_addr; // @[TensorStore.scala 152:16:@23954.4]
  wire [63:0] tensorFile_0_1__T_836_data; // @[TensorStore.scala 152:16:@23954.4]
  wire [10:0] tensorFile_0_1__T_836_addr; // @[TensorStore.scala 152:16:@23954.4]
  wire  tensorFile_0_1__T_836_mask; // @[TensorStore.scala 152:16:@23954.4]
  wire  tensorFile_0_1__T_836_en; // @[TensorStore.scala 152:16:@23954.4]
  wire [15:0] dec_sram_offset; // @[TensorStore.scala 51:29:@23729.4]
  wire [31:0] dec_dram_offset; // @[TensorStore.scala 51:29:@23731.4]
  wire [15:0] dec_ysize; // @[TensorStore.scala 51:29:@23735.4]
  wire [15:0] dec_xsize; // @[TensorStore.scala 51:29:@23737.4]
  wire [15:0] dec_xstride; // @[TensorStore.scala 51:29:@23739.4]
  reg [31:0] waddr_cur; // @[TensorStore.scala 52:22:@23749.4]
  reg [31:0] _RAND_2;
  reg [31:0] waddr_nxt; // @[TensorStore.scala 53:22:@23750.4]
  reg [31:0] _RAND_3;
  reg [7:0] xcnt; // @[TensorStore.scala 54:17:@23751.4]
  reg [31:0] _RAND_4;
  reg [7:0] xlen; // @[TensorStore.scala 55:17:@23752.4]
  reg [31:0] _RAND_5;
  reg [15:0] xrem; // @[TensorStore.scala 56:17:@23753.4]
  reg [31:0] _RAND_6;
  wire [16:0] _GEN_96; // @[TensorStore.scala 57:26:@23754.4]
  wire [16:0] _T_610; // @[TensorStore.scala 57:26:@23754.4]
  wire [17:0] _T_612; // @[TensorStore.scala 57:67:@23755.4]
  wire [17:0] _T_613; // @[TensorStore.scala 57:67:@23756.4]
  wire [16:0] xsize; // @[TensorStore.scala 57:67:@23757.4]
  reg [15:0] ycnt; // @[TensorStore.scala 60:17:@23758.4]
  reg [31:0] _RAND_7;
  reg [7:0] tag; // @[TensorStore.scala 62:16:@23759.4]
  reg [31:0] _RAND_8;
  reg [7:0] set; // @[TensorStore.scala 63:16:@23760.4]
  reg [31:0] _RAND_9;
  reg [31:0] xfer_bytes; // @[TensorStore.scala 65:23:@23761.4]
  reg [31:0] _RAND_10;
  wire [19:0] _GEN_97; // @[TensorStore.scala 66:35:@23762.4]
  wire [19:0] xstride_bytes; // @[TensorStore.scala 66:35:@23762.4]
  wire [35:0] _GEN_98; // @[TensorStore.scala 71:66:@23827.4]
  wire [35:0] _T_718; // @[TensorStore.scala 71:66:@23827.4]
  wire [35:0] _T_719; // @[TensorStore.scala 71:47:@23828.4]
  wire [35:0] _GEN_99; // @[TensorStore.scala 71:33:@23829.4]
  wire [35:0] xfer_init_addr; // @[TensorStore.scala 71:33:@23829.4]
  wire [32:0] _T_720; // @[TensorStore.scala 72:35:@23830.4]
  wire [31:0] xfer_split_addr; // @[TensorStore.scala 72:35:@23831.4]
  wire [31:0] _GEN_100; // @[TensorStore.scala 73:36:@23832.4]
  wire [32:0] _T_721; // @[TensorStore.scala 73:36:@23832.4]
  wire [31:0] xfer_stride_addr; // @[TensorStore.scala 73:36:@23833.4]
  wire [35:0] _GEN_15; // @[TensorStore.scala 75:55:@23834.4]
  wire [11:0] _T_722; // @[TensorStore.scala 75:55:@23834.4]
  wire [12:0] _T_723; // @[TensorStore.scala 75:38:@23835.4]
  wire [12:0] _T_724; // @[TensorStore.scala 75:38:@23836.4]
  wire [11:0] xfer_init_bytes; // @[TensorStore.scala 75:38:@23837.4]
  wire [8:0] xfer_init_pulses; // @[TensorStore.scala 76:43:@23838.4]
  wire [31:0] _GEN_16; // @[TensorStore.scala 77:56:@23839.4]
  wire [11:0] _T_725; // @[TensorStore.scala 77:56:@23839.4]
  wire [12:0] _T_726; // @[TensorStore.scala 77:38:@23840.4]
  wire [12:0] _T_727; // @[TensorStore.scala 77:38:@23841.4]
  wire [11:0] xfer_split_bytes; // @[TensorStore.scala 77:38:@23842.4]
  wire [8:0] xfer_split_pulses; // @[TensorStore.scala 78:44:@23843.4]
  wire [31:0] _GEN_43; // @[TensorStore.scala 79:57:@23844.4]
  wire [11:0] _T_728; // @[TensorStore.scala 79:57:@23844.4]
  wire [12:0] _T_729; // @[TensorStore.scala 79:38:@23845.4]
  wire [12:0] _T_730; // @[TensorStore.scala 79:38:@23846.4]
  wire [11:0] xfer_stride_bytes; // @[TensorStore.scala 79:38:@23847.4]
  wire [8:0] xfer_stride_pulses; // @[TensorStore.scala 80:45:@23848.4]
  reg [2:0] state; // @[TensorStore.scala 83:22:@23849.4]
  reg [31:0] _RAND_11;
  wire  _T_732; // @[Conditional.scala 37:30:@23850.4]
  wire [16:0] _GEN_101; // @[TensorStore.scala 91:21:@23855.8]
  wire  _T_733; // @[TensorStore.scala 91:21:@23855.8]
  wire [9:0] _T_736; // @[TensorStore.scala 95:36:@23861.10]
  wire [9:0] _T_737; // @[TensorStore.scala 95:36:@23862.10]
  wire [8:0] _T_738; // @[TensorStore.scala 95:36:@23863.10]
  wire [17:0] _T_739; // @[TensorStore.scala 96:25:@23865.10]
  wire [17:0] _T_740; // @[TensorStore.scala 96:25:@23866.10]
  wire [16:0] _T_741; // @[TensorStore.scala 96:25:@23867.10]
  wire [16:0] _GEN_0; // @[TensorStore.scala 91:41:@23856.8]
  wire [16:0] _GEN_1; // @[TensorStore.scala 91:41:@23856.8]
  wire [2:0] _GEN_2; // @[TensorStore.scala 89:23:@23853.6]
  wire [16:0] _GEN_3; // @[TensorStore.scala 89:23:@23853.6]
  wire [16:0] _GEN_4; // @[TensorStore.scala 89:23:@23853.6]
  wire  _T_742; // @[Conditional.scala 37:30:@23873.6]
  wire [2:0] _GEN_5; // @[TensorStore.scala 101:33:@23875.8]
  wire  _T_743; // @[Conditional.scala 37:30:@23880.8]
  wire  _T_744; // @[TensorStore.scala 107:19:@23883.12]
  wire  _T_746; // @[TensorStore.scala 109:24:@23888.14]
  wire [2:0] _GEN_6; // @[TensorStore.scala 109:49:@23889.14]
  wire [2:0] _GEN_7; // @[TensorStore.scala 107:29:@23884.12]
  wire [2:0] _GEN_8; // @[TensorStore.scala 106:34:@23882.10]
  wire  _T_747; // @[Conditional.scala 37:30:@23895.10]
  wire  _T_748; // @[Conditional.scala 37:30:@23900.12]
  wire  _T_750; // @[TensorStore.scala 119:19:@23903.16]
  wire [16:0] _T_752; // @[TensorStore.scala 120:31:@23905.18]
  wire [16:0] _T_753; // @[TensorStore.scala 120:31:@23906.18]
  wire [15:0] _T_754; // @[TensorStore.scala 120:31:@23907.18]
  wire  _T_755; // @[TensorStore.scala 120:21:@23908.18]
  wire [16:0] _GEN_103; // @[TensorStore.scala 125:24:@23915.20]
  wire  _T_756; // @[TensorStore.scala 125:24:@23915.20]
  wire [9:0] _T_759; // @[TensorStore.scala 129:42:@23921.22]
  wire [9:0] _T_760; // @[TensorStore.scala 129:42:@23922.22]
  wire [8:0] _T_761; // @[TensorStore.scala 129:42:@23923.22]
  wire [17:0] _T_762; // @[TensorStore.scala 130:29:@23925.22]
  wire [17:0] _T_763; // @[TensorStore.scala 130:29:@23926.22]
  wire [16:0] _T_764; // @[TensorStore.scala 130:29:@23927.22]
  wire [16:0] _GEN_9; // @[TensorStore.scala 125:46:@23916.20]
  wire [16:0] _GEN_10; // @[TensorStore.scala 125:46:@23916.20]
  wire [2:0] _GEN_11; // @[TensorStore.scala 120:38:@23909.18]
  wire [31:0] _GEN_12; // @[TensorStore.scala 120:38:@23909.18]
  wire [16:0] _GEN_13; // @[TensorStore.scala 120:38:@23909.18]
  wire [16:0] _GEN_14; // @[TensorStore.scala 120:38:@23909.18]
  wire [15:0] _GEN_105; // @[TensorStore.scala 134:24:@23933.18]
  wire  _T_765; // @[TensorStore.scala 134:24:@23933.18]
  wire [9:0] _T_768; // @[TensorStore.scala 143:37:@23943.20]
  wire [9:0] _T_769; // @[TensorStore.scala 143:37:@23944.20]
  wire [8:0] _T_770; // @[TensorStore.scala 143:37:@23945.20]
  wire [16:0] _T_771; // @[TensorStore.scala 144:24:@23947.20]
  wire [16:0] _T_772; // @[TensorStore.scala 144:24:@23948.20]
  wire [15:0] _T_773; // @[TensorStore.scala 144:24:@23949.20]
  wire [15:0] _GEN_17; // @[TensorStore.scala 134:45:@23934.18]
  wire [15:0] _GEN_18; // @[TensorStore.scala 134:45:@23934.18]
  wire [2:0] _GEN_19; // @[TensorStore.scala 119:28:@23904.16]
  wire [31:0] _GEN_20; // @[TensorStore.scala 119:28:@23904.16]
  wire [16:0] _GEN_21; // @[TensorStore.scala 119:28:@23904.16]
  wire [16:0] _GEN_22; // @[TensorStore.scala 119:28:@23904.16]
  wire [2:0] _GEN_23; // @[TensorStore.scala 118:27:@23902.14]
  wire [31:0] _GEN_24; // @[TensorStore.scala 118:27:@23902.14]
  wire [16:0] _GEN_25; // @[TensorStore.scala 118:27:@23902.14]
  wire [16:0] _GEN_26; // @[TensorStore.scala 118:27:@23902.14]
  wire [2:0] _GEN_27; // @[Conditional.scala 39:67:@23901.12]
  wire [31:0] _GEN_28; // @[Conditional.scala 39:67:@23901.12]
  wire [16:0] _GEN_29; // @[Conditional.scala 39:67:@23901.12]
  wire [16:0] _GEN_30; // @[Conditional.scala 39:67:@23901.12]
  wire [2:0] _GEN_31; // @[Conditional.scala 39:67:@23896.10]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67:@23896.10]
  wire [16:0] _GEN_33; // @[Conditional.scala 39:67:@23896.10]
  wire [16:0] _GEN_34; // @[Conditional.scala 39:67:@23896.10]
  wire [2:0] _GEN_35; // @[Conditional.scala 39:67:@23881.8]
  wire [31:0] _GEN_36; // @[Conditional.scala 39:67:@23881.8]
  wire [16:0] _GEN_37; // @[Conditional.scala 39:67:@23881.8]
  wire [16:0] _GEN_38; // @[Conditional.scala 39:67:@23881.8]
  wire [2:0] _GEN_39; // @[Conditional.scala 39:67:@23874.6]
  wire [31:0] _GEN_40; // @[Conditional.scala 39:67:@23874.6]
  wire [16:0] _GEN_41; // @[Conditional.scala 39:67:@23874.6]
  wire [16:0] _GEN_42; // @[Conditional.scala 39:67:@23874.6]
  wire [2:0] _GEN_44; // @[Conditional.scala 40:58:@23851.4]
  wire [16:0] _GEN_45; // @[Conditional.scala 40:58:@23851.4]
  wire [16:0] _GEN_46; // @[Conditional.scala 40:58:@23851.4]
  wire [63:0] _T_804; // @[TensorStore.scala 163:46:@23967.4]
  wire [127:0] _T_812; // @[TensorStore.scala 163:46:@23975.4]
  wire  _T_844; // @[TensorStore.scala 170:22:@23992.4]
  wire  _T_845; // @[TensorStore.scala 170:36:@23993.4]
  wire [8:0] _T_847; // @[TensorStore.scala 172:19:@23994.4]
  wire [7:0] _T_848; // @[TensorStore.scala 172:19:@23995.4]
  wire  _T_849; // @[TensorStore.scala 172:10:@23996.4]
  wire  _T_850; // @[TensorStore.scala 171:19:@23997.4]
  wire  _T_853; // @[TensorStore.scala 172:25:@23999.4]
  wire  _T_858; // @[TensorStore.scala 174:10:@24003.4]
  wire  stride; // @[TensorStore.scala 173:18:@24004.4]
  wire  _T_859; // @[TensorStore.scala 176:14:@24005.4]
  wire [16:0] _T_862; // @[TensorStore.scala 179:18:@24011.8]
  wire [15:0] _T_863; // @[TensorStore.scala 179:18:@24012.8]
  wire [15:0] _GEN_58; // @[TensorStore.scala 178:22:@24010.6]
  wire  _T_864; // @[TensorStore.scala 182:14:@24015.4]
  wire  _T_867; // @[TensorStore.scala 182:28:@24017.4]
  wire  _T_869; // @[Decoupled.scala 37:37:@24022.6]
  wire [8:0] _T_871; // @[TensorStore.scala 185:16:@24024.8]
  wire [7:0] _T_872; // @[TensorStore.scala 185:16:@24025.8]
  wire [7:0] _GEN_60; // @[TensorStore.scala 184:37:@24023.6]
  wire  _T_875; // @[TensorStore.scala 189:33:@24029.4]
  wire  _T_878; // @[TensorStore.scala 189:58:@24031.4]
  wire  _T_879; // @[TensorStore.scala 189:25:@24032.4]
  wire  _T_884; // @[TensorStore.scala 191:36:@24039.6]
  wire [8:0] _T_886; // @[TensorStore.scala 192:16:@24041.8]
  wire [7:0] _T_887; // @[TensorStore.scala 192:16:@24042.8]
  wire [7:0] _GEN_62; // @[TensorStore.scala 191:68:@24040.6]
  reg [10:0] raddr_cur; // @[TensorStore.scala 195:22:@24045.4]
  reg [31:0] _RAND_12;
  reg [10:0] raddr_nxt; // @[TensorStore.scala 196:22:@24046.4]
  reg [31:0] _RAND_13;
  wire  _T_894; // @[TensorStore.scala 200:36:@24055.6]
  wire  _T_897; // @[TensorStore.scala 200:68:@24057.6]
  wire [11:0] _T_899; // @[TensorStore.scala 201:28:@24059.8]
  wire [10:0] _T_900; // @[TensorStore.scala 201:28:@24060.8]
  wire [15:0] _GEN_107; // @[TensorStore.scala 203:28:@24065.10]
  wire [16:0] _T_901; // @[TensorStore.scala 203:28:@24065.10]
  wire [15:0] _T_902; // @[TensorStore.scala 203:28:@24066.10]
  wire [15:0] _GEN_64; // @[TensorStore.scala 202:22:@24064.8]
  wire [15:0] _GEN_65; // @[TensorStore.scala 202:22:@24064.8]
  wire [15:0] _GEN_66; // @[TensorStore.scala 200:100:@24058.6]
  wire [15:0] _GEN_67; // @[TensorStore.scala 200:100:@24058.6]
  wire [15:0] _GEN_68; // @[TensorStore.scala 197:25:@24048.4]
  wire [15:0] _GEN_69; // @[TensorStore.scala 197:25:@24048.4]
  wire  _T_907; // @[TensorStore.scala 209:65:@24073.4]
  wire  _T_908; // @[TensorStore.scala 209:57:@24074.4]
  wire  _GEN_71; // @[TensorStore.scala 209:25:@24077.4]
  wire  _T_960; // @[Mux.scala 46:19:@24090.4]
  wire [63:0] mdata_0; // @[Mux.scala 46:16:@24091.4]
  wire [63:0] mdata_1; // @[Mux.scala 46:16:@24091.4]
  wire  _T_975; // @[TensorStore.scala 217:59:@24100.6]
  wire  _T_976; // @[TensorStore.scala 217:51:@24101.6]
  wire [31:0] _GEN_74; // @[TensorStore.scala 219:22:@24106.8]
  wire [31:0] _GEN_75; // @[TensorStore.scala 219:22:@24106.8]
  wire [31:0] _GEN_76; // @[TensorStore.scala 217:68:@24102.6]
  wire [31:0] _GEN_77; // @[TensorStore.scala 217:68:@24102.6]
  wire [35:0] _GEN_78; // @[TensorStore.scala 214:25:@24093.4]
  wire [35:0] _GEN_79; // @[TensorStore.scala 214:25:@24093.4]
  wire  _T_982; // @[:@24116.4]
  wire [8:0] _T_987; // @[TensorStore.scala 234:18:@24125.8]
  wire [7:0] _T_988; // @[TensorStore.scala 234:18:@24126.8]
  wire [7:0] _GEN_82; // @[TensorStore.scala 233:37:@24124.6]
  wire  _T_1010; // @[TensorStore.scala 241:50:@24149.4]
  reg [10:0] tensorFile_0_0__T_914_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [10:0] tensorFile_0_1__T_914_addr_pipe_0;
  reg [31:0] _RAND_15;
  assign tensorFile_0_0__T_914_addr = tensorFile_0_0__T_914_addr_pipe_0;
  assign tensorFile_0_0__T_914_data = tensorFile_0_0[tensorFile_0_0__T_914_addr]; // @[TensorStore.scala 152:16:@23954.4]
  assign tensorFile_0_0__T_836_data = _T_812[63:0];
  assign tensorFile_0_0__T_836_addr = io_tensor_wr_bits_idx;
  assign tensorFile_0_0__T_836_mask = 1'h1;
  assign tensorFile_0_0__T_836_en = io_tensor_wr_valid;
  assign tensorFile_0_1__T_914_addr = tensorFile_0_1__T_914_addr_pipe_0;
  assign tensorFile_0_1__T_914_data = tensorFile_0_1[tensorFile_0_1__T_914_addr]; // @[TensorStore.scala 152:16:@23954.4]
  assign tensorFile_0_1__T_836_data = _T_812[127:64];
  assign tensorFile_0_1__T_836_addr = io_tensor_wr_bits_idx;
  assign tensorFile_0_1__T_836_mask = 1'h1;
  assign tensorFile_0_1__T_836_en = io_tensor_wr_valid;
  assign dec_sram_offset = io_inst[24:9]; // @[TensorStore.scala 51:29:@23729.4]
  assign dec_dram_offset = io_inst[56:25]; // @[TensorStore.scala 51:29:@23731.4]
  assign dec_ysize = io_inst[79:64]; // @[TensorStore.scala 51:29:@23735.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorStore.scala 51:29:@23737.4]
  assign dec_xstride = io_inst[111:96]; // @[TensorStore.scala 51:29:@23739.4]
  assign _GEN_96 = {{1'd0}, dec_xsize}; // @[TensorStore.scala 57:26:@23754.4]
  assign _T_610 = _GEN_96 << 1; // @[TensorStore.scala 57:26:@23754.4]
  assign _T_612 = _T_610 - 17'h1; // @[TensorStore.scala 57:67:@23755.4]
  assign _T_613 = $unsigned(_T_612); // @[TensorStore.scala 57:67:@23756.4]
  assign xsize = _T_613[16:0]; // @[TensorStore.scala 57:67:@23757.4]
  assign _GEN_97 = {{4'd0}, dec_xstride}; // @[TensorStore.scala 66:35:@23762.4]
  assign xstride_bytes = _GEN_97 << 4; // @[TensorStore.scala 66:35:@23762.4]
  assign _GEN_98 = {{4'd0}, dec_dram_offset}; // @[TensorStore.scala 71:66:@23827.4]
  assign _T_718 = _GEN_98 << 4; // @[TensorStore.scala 71:66:@23827.4]
  assign _T_719 = 36'hffffffff & _T_718; // @[TensorStore.scala 71:47:@23828.4]
  assign _GEN_99 = {{4'd0}, io_baddr}; // @[TensorStore.scala 71:33:@23829.4]
  assign xfer_init_addr = _GEN_99 | _T_719; // @[TensorStore.scala 71:33:@23829.4]
  assign _T_720 = waddr_cur + xfer_bytes; // @[TensorStore.scala 72:35:@23830.4]
  assign xfer_split_addr = waddr_cur + xfer_bytes; // @[TensorStore.scala 72:35:@23831.4]
  assign _GEN_100 = {{12'd0}, xstride_bytes}; // @[TensorStore.scala 73:36:@23832.4]
  assign _T_721 = waddr_nxt + _GEN_100; // @[TensorStore.scala 73:36:@23832.4]
  assign xfer_stride_addr = waddr_nxt + _GEN_100; // @[TensorStore.scala 73:36:@23833.4]
  assign _GEN_15 = xfer_init_addr % 36'h800; // @[TensorStore.scala 75:55:@23834.4]
  assign _T_722 = _GEN_15[11:0]; // @[TensorStore.scala 75:55:@23834.4]
  assign _T_723 = 12'h800 - _T_722; // @[TensorStore.scala 75:38:@23835.4]
  assign _T_724 = $unsigned(_T_723); // @[TensorStore.scala 75:38:@23836.4]
  assign xfer_init_bytes = _T_724[11:0]; // @[TensorStore.scala 75:38:@23837.4]
  assign xfer_init_pulses = xfer_init_bytes[11:3]; // @[TensorStore.scala 76:43:@23838.4]
  assign _GEN_16 = xfer_split_addr % 32'h800; // @[TensorStore.scala 77:56:@23839.4]
  assign _T_725 = _GEN_16[11:0]; // @[TensorStore.scala 77:56:@23839.4]
  assign _T_726 = 12'h800 - _T_725; // @[TensorStore.scala 77:38:@23840.4]
  assign _T_727 = $unsigned(_T_726); // @[TensorStore.scala 77:38:@23841.4]
  assign xfer_split_bytes = _T_727[11:0]; // @[TensorStore.scala 77:38:@23842.4]
  assign xfer_split_pulses = xfer_split_bytes[11:3]; // @[TensorStore.scala 78:44:@23843.4]
  assign _GEN_43 = xfer_stride_addr % 32'h800; // @[TensorStore.scala 79:57:@23844.4]
  assign _T_728 = _GEN_43[11:0]; // @[TensorStore.scala 79:57:@23844.4]
  assign _T_729 = 12'h800 - _T_728; // @[TensorStore.scala 79:38:@23845.4]
  assign _T_730 = $unsigned(_T_729); // @[TensorStore.scala 79:38:@23846.4]
  assign xfer_stride_bytes = _T_730[11:0]; // @[TensorStore.scala 79:38:@23847.4]
  assign xfer_stride_pulses = xfer_stride_bytes[11:3]; // @[TensorStore.scala 80:45:@23848.4]
  assign _T_732 = 3'h0 == state; // @[Conditional.scala 37:30:@23850.4]
  assign _GEN_101 = {{8'd0}, xfer_init_pulses}; // @[TensorStore.scala 91:21:@23855.8]
  assign _T_733 = xsize < _GEN_101; // @[TensorStore.scala 91:21:@23855.8]
  assign _T_736 = xfer_init_pulses - 9'h1; // @[TensorStore.scala 95:36:@23861.10]
  assign _T_737 = $unsigned(_T_736); // @[TensorStore.scala 95:36:@23862.10]
  assign _T_738 = _T_737[8:0]; // @[TensorStore.scala 95:36:@23863.10]
  assign _T_739 = xsize - _GEN_101; // @[TensorStore.scala 96:25:@23865.10]
  assign _T_740 = $unsigned(_T_739); // @[TensorStore.scala 96:25:@23866.10]
  assign _T_741 = _T_740[16:0]; // @[TensorStore.scala 96:25:@23867.10]
  assign _GEN_0 = _T_733 ? xsize : {{8'd0}, _T_738}; // @[TensorStore.scala 91:41:@23856.8]
  assign _GEN_1 = _T_733 ? 17'h0 : _T_741; // @[TensorStore.scala 91:41:@23856.8]
  assign _GEN_2 = io_start ? 3'h1 : state; // @[TensorStore.scala 89:23:@23853.6]
  assign _GEN_3 = io_start ? _GEN_0 : {{9'd0}, xlen}; // @[TensorStore.scala 89:23:@23853.6]
  assign _GEN_4 = io_start ? _GEN_1 : {{1'd0}, xrem}; // @[TensorStore.scala 89:23:@23853.6]
  assign _T_742 = 3'h1 == state; // @[Conditional.scala 37:30:@23873.6]
  assign _GEN_5 = io_vme_wr_cmd_ready ? 3'h2 : state; // @[TensorStore.scala 101:33:@23875.8]
  assign _T_743 = 3'h2 == state; // @[Conditional.scala 37:30:@23880.8]
  assign _T_744 = xcnt == xlen; // @[TensorStore.scala 107:19:@23883.12]
  assign _T_746 = tag == 8'h1; // @[TensorStore.scala 109:24:@23888.14]
  assign _GEN_6 = _T_746 ? 3'h3 : state; // @[TensorStore.scala 109:49:@23889.14]
  assign _GEN_7 = _T_744 ? 3'h4 : _GEN_6; // @[TensorStore.scala 107:29:@23884.12]
  assign _GEN_8 = io_vme_wr_data_ready ? _GEN_7 : state; // @[TensorStore.scala 106:34:@23882.10]
  assign _T_747 = 3'h3 == state; // @[Conditional.scala 37:30:@23895.10]
  assign _T_748 = 3'h4 == state; // @[Conditional.scala 37:30:@23900.12]
  assign _T_750 = xrem == 16'h0; // @[TensorStore.scala 119:19:@23903.16]
  assign _T_752 = dec_ysize - 16'h1; // @[TensorStore.scala 120:31:@23905.18]
  assign _T_753 = $unsigned(_T_752); // @[TensorStore.scala 120:31:@23906.18]
  assign _T_754 = _T_753[15:0]; // @[TensorStore.scala 120:31:@23907.18]
  assign _T_755 = ycnt == _T_754; // @[TensorStore.scala 120:21:@23908.18]
  assign _GEN_103 = {{8'd0}, xfer_stride_pulses}; // @[TensorStore.scala 125:24:@23915.20]
  assign _T_756 = xsize < _GEN_103; // @[TensorStore.scala 125:24:@23915.20]
  assign _T_759 = xfer_stride_pulses - 9'h1; // @[TensorStore.scala 129:42:@23921.22]
  assign _T_760 = $unsigned(_T_759); // @[TensorStore.scala 129:42:@23922.22]
  assign _T_761 = _T_760[8:0]; // @[TensorStore.scala 129:42:@23923.22]
  assign _T_762 = xsize - _GEN_103; // @[TensorStore.scala 130:29:@23925.22]
  assign _T_763 = $unsigned(_T_762); // @[TensorStore.scala 130:29:@23926.22]
  assign _T_764 = _T_763[16:0]; // @[TensorStore.scala 130:29:@23927.22]
  assign _GEN_9 = _T_756 ? xsize : {{8'd0}, _T_761}; // @[TensorStore.scala 125:46:@23916.20]
  assign _GEN_10 = _T_756 ? 17'h0 : _T_764; // @[TensorStore.scala 125:46:@23916.20]
  assign _GEN_11 = _T_755 ? 3'h0 : 3'h1; // @[TensorStore.scala 120:38:@23909.18]
  assign _GEN_12 = _T_755 ? xfer_bytes : {{20'd0}, xfer_stride_bytes}; // @[TensorStore.scala 120:38:@23909.18]
  assign _GEN_13 = _T_755 ? {{9'd0}, xlen} : _GEN_9; // @[TensorStore.scala 120:38:@23909.18]
  assign _GEN_14 = _T_755 ? {{1'd0}, xrem} : _GEN_10; // @[TensorStore.scala 120:38:@23909.18]
  assign _GEN_105 = {{7'd0}, xfer_split_pulses}; // @[TensorStore.scala 134:24:@23933.18]
  assign _T_765 = xrem < _GEN_105; // @[TensorStore.scala 134:24:@23933.18]
  assign _T_768 = xfer_split_pulses - 9'h1; // @[TensorStore.scala 143:37:@23943.20]
  assign _T_769 = $unsigned(_T_768); // @[TensorStore.scala 143:37:@23944.20]
  assign _T_770 = _T_769[8:0]; // @[TensorStore.scala 143:37:@23945.20]
  assign _T_771 = xrem - _GEN_105; // @[TensorStore.scala 144:24:@23947.20]
  assign _T_772 = $unsigned(_T_771); // @[TensorStore.scala 144:24:@23948.20]
  assign _T_773 = _T_772[15:0]; // @[TensorStore.scala 144:24:@23949.20]
  assign _GEN_17 = _T_765 ? xrem : {{7'd0}, _T_770}; // @[TensorStore.scala 134:45:@23934.18]
  assign _GEN_18 = _T_765 ? 16'h0 : _T_773; // @[TensorStore.scala 134:45:@23934.18]
  assign _GEN_19 = _T_750 ? _GEN_11 : 3'h1; // @[TensorStore.scala 119:28:@23904.16]
  assign _GEN_20 = _T_750 ? _GEN_12 : {{20'd0}, xfer_split_bytes}; // @[TensorStore.scala 119:28:@23904.16]
  assign _GEN_21 = _T_750 ? _GEN_13 : {{1'd0}, _GEN_17}; // @[TensorStore.scala 119:28:@23904.16]
  assign _GEN_22 = _T_750 ? _GEN_14 : {{1'd0}, _GEN_18}; // @[TensorStore.scala 119:28:@23904.16]
  assign _GEN_23 = io_vme_wr_ack ? _GEN_19 : state; // @[TensorStore.scala 118:27:@23902.14]
  assign _GEN_24 = io_vme_wr_ack ? _GEN_20 : xfer_bytes; // @[TensorStore.scala 118:27:@23902.14]
  assign _GEN_25 = io_vme_wr_ack ? _GEN_21 : {{9'd0}, xlen}; // @[TensorStore.scala 118:27:@23902.14]
  assign _GEN_26 = io_vme_wr_ack ? _GEN_22 : {{1'd0}, xrem}; // @[TensorStore.scala 118:27:@23902.14]
  assign _GEN_27 = _T_748 ? _GEN_23 : state; // @[Conditional.scala 39:67:@23901.12]
  assign _GEN_28 = _T_748 ? _GEN_24 : xfer_bytes; // @[Conditional.scala 39:67:@23901.12]
  assign _GEN_29 = _T_748 ? _GEN_25 : {{9'd0}, xlen}; // @[Conditional.scala 39:67:@23901.12]
  assign _GEN_30 = _T_748 ? _GEN_26 : {{1'd0}, xrem}; // @[Conditional.scala 39:67:@23901.12]
  assign _GEN_31 = _T_747 ? 3'h2 : _GEN_27; // @[Conditional.scala 39:67:@23896.10]
  assign _GEN_32 = _T_747 ? xfer_bytes : _GEN_28; // @[Conditional.scala 39:67:@23896.10]
  assign _GEN_33 = _T_747 ? {{9'd0}, xlen} : _GEN_29; // @[Conditional.scala 39:67:@23896.10]
  assign _GEN_34 = _T_747 ? {{1'd0}, xrem} : _GEN_30; // @[Conditional.scala 39:67:@23896.10]
  assign _GEN_35 = _T_743 ? _GEN_8 : _GEN_31; // @[Conditional.scala 39:67:@23881.8]
  assign _GEN_36 = _T_743 ? xfer_bytes : _GEN_32; // @[Conditional.scala 39:67:@23881.8]
  assign _GEN_37 = _T_743 ? {{9'd0}, xlen} : _GEN_33; // @[Conditional.scala 39:67:@23881.8]
  assign _GEN_38 = _T_743 ? {{1'd0}, xrem} : _GEN_34; // @[Conditional.scala 39:67:@23881.8]
  assign _GEN_39 = _T_742 ? _GEN_5 : _GEN_35; // @[Conditional.scala 39:67:@23874.6]
  assign _GEN_40 = _T_742 ? xfer_bytes : _GEN_36; // @[Conditional.scala 39:67:@23874.6]
  assign _GEN_41 = _T_742 ? {{9'd0}, xlen} : _GEN_37; // @[Conditional.scala 39:67:@23874.6]
  assign _GEN_42 = _T_742 ? {{1'd0}, xrem} : _GEN_38; // @[Conditional.scala 39:67:@23874.6]
  assign _GEN_44 = _T_732 ? _GEN_2 : _GEN_39; // @[Conditional.scala 40:58:@23851.4]
  assign _GEN_45 = _T_732 ? _GEN_3 : _GEN_41; // @[Conditional.scala 40:58:@23851.4]
  assign _GEN_46 = _T_732 ? _GEN_4 : _GEN_42; // @[Conditional.scala 40:58:@23851.4]
  assign _T_804 = {io_tensor_wr_bits_data_0_7,io_tensor_wr_bits_data_0_6,io_tensor_wr_bits_data_0_5,io_tensor_wr_bits_data_0_4,io_tensor_wr_bits_data_0_3,io_tensor_wr_bits_data_0_2,io_tensor_wr_bits_data_0_1,io_tensor_wr_bits_data_0_0}; // @[TensorStore.scala 163:46:@23967.4]
  assign _T_812 = {io_tensor_wr_bits_data_0_15,io_tensor_wr_bits_data_0_14,io_tensor_wr_bits_data_0_13,io_tensor_wr_bits_data_0_12,io_tensor_wr_bits_data_0_11,io_tensor_wr_bits_data_0_10,io_tensor_wr_bits_data_0_9,io_tensor_wr_bits_data_0_8,_T_804}; // @[TensorStore.scala 163:46:@23975.4]
  assign _T_844 = state == 3'h4; // @[TensorStore.scala 170:22:@23992.4]
  assign _T_845 = _T_844 & io_vme_wr_ack; // @[TensorStore.scala 170:36:@23993.4]
  assign _T_847 = xlen + 8'h1; // @[TensorStore.scala 172:19:@23994.4]
  assign _T_848 = xlen + 8'h1; // @[TensorStore.scala 172:19:@23995.4]
  assign _T_849 = xcnt == _T_848; // @[TensorStore.scala 172:10:@23996.4]
  assign _T_850 = _T_845 & _T_849; // @[TensorStore.scala 171:19:@23997.4]
  assign _T_853 = _T_850 & _T_750; // @[TensorStore.scala 172:25:@23999.4]
  assign _T_858 = ycnt != _T_754; // @[TensorStore.scala 174:10:@24003.4]
  assign stride = _T_853 & _T_858; // @[TensorStore.scala 173:18:@24004.4]
  assign _T_859 = state == 3'h0; // @[TensorStore.scala 176:14:@24005.4]
  assign _T_862 = ycnt + 16'h1; // @[TensorStore.scala 179:18:@24011.8]
  assign _T_863 = ycnt + 16'h1; // @[TensorStore.scala 179:18:@24012.8]
  assign _GEN_58 = stride ? _T_863 : ycnt; // @[TensorStore.scala 178:22:@24010.6]
  assign _T_864 = state == 3'h1; // @[TensorStore.scala 182:14:@24015.4]
  assign _T_867 = _T_864 | _T_746; // @[TensorStore.scala 182:28:@24017.4]
  assign _T_869 = io_vme_wr_data_ready & io_vme_wr_data_valid; // @[Decoupled.scala 37:37:@24022.6]
  assign _T_871 = tag + 8'h1; // @[TensorStore.scala 185:16:@24024.8]
  assign _T_872 = tag + 8'h1; // @[TensorStore.scala 185:16:@24025.8]
  assign _GEN_60 = _T_869 ? _T_872 : tag; // @[TensorStore.scala 184:37:@24023.6]
  assign _T_875 = set == 8'h0; // @[TensorStore.scala 189:33:@24029.4]
  assign _T_878 = _T_875 & _T_746; // @[TensorStore.scala 189:58:@24031.4]
  assign _T_879 = _T_864 | _T_878; // @[TensorStore.scala 189:25:@24032.4]
  assign _T_884 = _T_869 & _T_746; // @[TensorStore.scala 191:36:@24039.6]
  assign _T_886 = set + 8'h1; // @[TensorStore.scala 192:16:@24041.8]
  assign _T_887 = set + 8'h1; // @[TensorStore.scala 192:16:@24042.8]
  assign _GEN_62 = _T_884 ? _T_887 : set; // @[TensorStore.scala 191:68:@24040.6]
  assign _T_894 = _T_869 & _T_875; // @[TensorStore.scala 200:36:@24055.6]
  assign _T_897 = _T_894 & _T_746; // @[TensorStore.scala 200:68:@24057.6]
  assign _T_899 = raddr_cur + 11'h1; // @[TensorStore.scala 201:28:@24059.8]
  assign _T_900 = raddr_cur + 11'h1; // @[TensorStore.scala 201:28:@24060.8]
  assign _GEN_107 = {{5'd0}, raddr_nxt}; // @[TensorStore.scala 203:28:@24065.10]
  assign _T_901 = _GEN_107 + dec_xsize; // @[TensorStore.scala 203:28:@24065.10]
  assign _T_902 = _GEN_107 + dec_xsize; // @[TensorStore.scala 203:28:@24066.10]
  assign _GEN_64 = stride ? _T_902 : {{5'd0}, raddr_cur}; // @[TensorStore.scala 202:22:@24064.8]
  assign _GEN_65 = stride ? _T_902 : {{5'd0}, raddr_nxt}; // @[TensorStore.scala 202:22:@24064.8]
  assign _GEN_66 = _T_897 ? {{5'd0}, _T_900} : _GEN_64; // @[TensorStore.scala 200:100:@24058.6]
  assign _GEN_67 = _T_897 ? {{5'd0}, raddr_nxt} : _GEN_65; // @[TensorStore.scala 200:100:@24058.6]
  assign _GEN_68 = _T_859 ? dec_sram_offset : _GEN_66; // @[TensorStore.scala 197:25:@24048.4]
  assign _GEN_69 = _T_859 ? dec_sram_offset : _GEN_67; // @[TensorStore.scala 197:25:@24048.4]
  assign _T_907 = state == 3'h3; // @[TensorStore.scala 209:65:@24073.4]
  assign _T_908 = _T_864 | _T_907; // @[TensorStore.scala 209:57:@24074.4]
  assign _GEN_71 = _T_908; // @[TensorStore.scala 209:25:@24077.4]
  assign _T_960 = 8'h0 == set; // @[Mux.scala 46:19:@24090.4]
  assign mdata_0 = _T_960 ? tensorFile_0_0__T_914_data : 64'h0; // @[Mux.scala 46:16:@24091.4]
  assign mdata_1 = _T_960 ? tensorFile_0_1__T_914_data : 64'h0; // @[Mux.scala 46:16:@24091.4]
  assign _T_975 = xrem != 16'h0; // @[TensorStore.scala 217:59:@24100.6]
  assign _T_976 = _T_845 & _T_975; // @[TensorStore.scala 217:51:@24101.6]
  assign _GEN_74 = stride ? xfer_stride_addr : waddr_cur; // @[TensorStore.scala 219:22:@24106.8]
  assign _GEN_75 = stride ? xfer_stride_addr : waddr_nxt; // @[TensorStore.scala 219:22:@24106.8]
  assign _GEN_76 = _T_976 ? xfer_split_addr : _GEN_74; // @[TensorStore.scala 217:68:@24102.6]
  assign _GEN_77 = _T_976 ? waddr_nxt : _GEN_75; // @[TensorStore.scala 217:68:@24102.6]
  assign _GEN_78 = _T_859 ? xfer_init_addr : {{4'd0}, _GEN_76}; // @[TensorStore.scala 214:25:@24093.4]
  assign _GEN_79 = _T_859 ? xfer_init_addr : {{4'd0}, _GEN_77}; // @[TensorStore.scala 214:25:@24093.4]
  assign _T_982 = tag[0]; // @[:@24116.4]
  assign _T_987 = xcnt + 8'h1; // @[TensorStore.scala 234:18:@24125.8]
  assign _T_988 = xcnt + 8'h1; // @[TensorStore.scala 234:18:@24126.8]
  assign _GEN_82 = _T_869 ? _T_988 : xcnt; // @[TensorStore.scala 233:37:@24124.6]
  assign _T_1010 = _T_845 & _T_750; // @[TensorStore.scala 241:50:@24149.4]
  assign io_done = _T_1010 & _T_755; // @[TensorStore.scala 241:11:@24155.4]
  assign io_vme_wr_cmd_valid = state == 3'h1; // @[TensorStore.scala 224:23:@24111.4]
  assign io_vme_wr_cmd_bits_addr = waddr_cur; // @[TensorStore.scala 225:27:@24112.4]
  assign io_vme_wr_cmd_bits_len = xlen; // @[TensorStore.scala 226:26:@24113.4]
  assign io_vme_wr_data_valid = state == 3'h2; // @[TensorStore.scala 228:24:@24115.4]
  assign io_vme_wr_data_bits = _T_982 ? mdata_1 : mdata_0; // @[TensorStore.scala 229:23:@24117.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_0[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_1[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  waddr_cur = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  waddr_nxt = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xcnt = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  xlen = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  xrem = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ycnt = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tag = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  set = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  xfer_bytes = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  raddr_cur = _RAND_12[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  raddr_nxt = _RAND_13[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  tensorFile_0_0__T_914_addr_pipe_0 = _RAND_14[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  tensorFile_0_1__T_914_addr_pipe_0 = _RAND_15[10:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tensorFile_0_0__T_836_en & tensorFile_0_0__T_836_mask) begin
      tensorFile_0_0[tensorFile_0_0__T_836_addr] <= tensorFile_0_0__T_836_data; // @[TensorStore.scala 152:16:@23954.4]
    end
    if(tensorFile_0_1__T_836_en & tensorFile_0_1__T_836_mask) begin
      tensorFile_0_1[tensorFile_0_1__T_836_addr] <= tensorFile_0_1__T_836_data; // @[TensorStore.scala 152:16:@23954.4]
    end
    waddr_cur <= _GEN_78[31:0];
    waddr_nxt <= _GEN_79[31:0];
    if (_T_864) begin
      xcnt <= 8'h0;
    end else begin
      if (_T_869) begin
        xcnt <= _T_988;
      end
    end
    xlen <= _GEN_45[7:0];
    xrem <= _GEN_46[15:0];
    if (_T_859) begin
      ycnt <= 16'h0;
    end else begin
      if (stride) begin
        ycnt <= _T_863;
      end
    end
    if (_T_867) begin
      tag <= 8'h0;
    end else begin
      if (_T_869) begin
        tag <= _T_872;
      end
    end
    if (_T_879) begin
      set <= 8'h0;
    end else begin
      if (_T_884) begin
        set <= _T_887;
      end
    end
    if (_T_732) begin
      xfer_bytes <= {{20'd0}, xfer_init_bytes};
    end else begin
      if (!(_T_742)) begin
        if (!(_T_743)) begin
          if (!(_T_747)) begin
            if (_T_748) begin
              if (io_vme_wr_ack) begin
                if (_T_750) begin
                  if (!(_T_755)) begin
                    xfer_bytes <= {{20'd0}, xfer_stride_bytes};
                  end
                end else begin
                  xfer_bytes <= {{20'd0}, xfer_split_bytes};
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_732) begin
        if (io_start) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_742) begin
          if (io_vme_wr_cmd_ready) begin
            state <= 3'h2;
          end
        end else begin
          if (_T_743) begin
            if (io_vme_wr_data_ready) begin
              if (_T_744) begin
                state <= 3'h4;
              end else begin
                if (_T_746) begin
                  state <= 3'h3;
                end
              end
            end
          end else begin
            if (_T_747) begin
              state <= 3'h2;
            end else begin
              if (_T_748) begin
                if (io_vme_wr_ack) begin
                  if (_T_750) begin
                    if (_T_755) begin
                      state <= 3'h0;
                    end else begin
                      state <= 3'h1;
                    end
                  end else begin
                    state <= 3'h1;
                  end
                end
              end
            end
          end
        end
      end
    end
    raddr_cur <= _GEN_68[10:0];
    raddr_nxt <= _GEN_69[10:0];
    if (_GEN_71) begin
      tensorFile_0_0__T_914_addr_pipe_0 <= raddr_cur;
    end
    if (_GEN_71) begin
      tensorFile_0_1__T_914_addr_pipe_0 <= raddr_cur;
    end
  end
endmodule
module Store( // @[:@24157.2]
  input          clock, // @[:@24158.4]
  input          reset, // @[:@24159.4]
  input          io_i_post, // @[:@24160.4]
  output         io_o_post, // @[:@24160.4]
  output         io_inst_ready, // @[:@24160.4]
  input          io_inst_valid, // @[:@24160.4]
  input  [127:0] io_inst_bits, // @[:@24160.4]
  input  [31:0]  io_out_baddr, // @[:@24160.4]
  input          io_vme_wr_cmd_ready, // @[:@24160.4]
  output         io_vme_wr_cmd_valid, // @[:@24160.4]
  output [31:0]  io_vme_wr_cmd_bits_addr, // @[:@24160.4]
  output [7:0]   io_vme_wr_cmd_bits_len, // @[:@24160.4]
  input          io_vme_wr_data_ready, // @[:@24160.4]
  output         io_vme_wr_data_valid, // @[:@24160.4]
  output [63:0]  io_vme_wr_data_bits, // @[:@24160.4]
  input          io_vme_wr_ack, // @[:@24160.4]
  input          io_out_wr_valid, // @[:@24160.4]
  input  [10:0]  io_out_wr_bits_idx, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_0, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_1, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_2, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_3, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_4, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_5, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_6, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_7, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_8, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_9, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_10, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_11, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_12, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_13, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_14, // @[:@24160.4]
  input  [7:0]   io_out_wr_bits_data_0_15 // @[:@24160.4]
);
  wire  s_clock; // @[Store.scala 46:17:@24163.4]
  wire  s_reset; // @[Store.scala 46:17:@24163.4]
  wire  s_io_spost; // @[Store.scala 46:17:@24163.4]
  wire  s_io_swait; // @[Store.scala 46:17:@24163.4]
  wire  s_io_sready; // @[Store.scala 46:17:@24163.4]
  wire  inst_q_clock; // @[Store.scala 47:22:@24166.4]
  wire  inst_q_reset; // @[Store.scala 47:22:@24166.4]
  wire  inst_q_io_enq_ready; // @[Store.scala 47:22:@24166.4]
  wire  inst_q_io_enq_valid; // @[Store.scala 47:22:@24166.4]
  wire [127:0] inst_q_io_enq_bits; // @[Store.scala 47:22:@24166.4]
  wire  inst_q_io_deq_ready; // @[Store.scala 47:22:@24166.4]
  wire  inst_q_io_deq_valid; // @[Store.scala 47:22:@24166.4]
  wire [127:0] inst_q_io_deq_bits; // @[Store.scala 47:22:@24166.4]
  wire [127:0] dec_io_inst; // @[Store.scala 49:19:@24169.4]
  wire  dec_io_push_prev; // @[Store.scala 49:19:@24169.4]
  wire  dec_io_pop_prev; // @[Store.scala 49:19:@24169.4]
  wire  dec_io_isStore; // @[Store.scala 49:19:@24169.4]
  wire  dec_io_isSync; // @[Store.scala 49:19:@24169.4]
  wire  tensorStore_clock; // @[Store.scala 52:27:@24173.4]
  wire  tensorStore_reset; // @[Store.scala 52:27:@24173.4]
  wire  tensorStore_io_start; // @[Store.scala 52:27:@24173.4]
  wire  tensorStore_io_done; // @[Store.scala 52:27:@24173.4]
  wire [127:0] tensorStore_io_inst; // @[Store.scala 52:27:@24173.4]
  wire [31:0] tensorStore_io_baddr; // @[Store.scala 52:27:@24173.4]
  wire  tensorStore_io_vme_wr_cmd_ready; // @[Store.scala 52:27:@24173.4]
  wire  tensorStore_io_vme_wr_cmd_valid; // @[Store.scala 52:27:@24173.4]
  wire [31:0] tensorStore_io_vme_wr_cmd_bits_addr; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_vme_wr_cmd_bits_len; // @[Store.scala 52:27:@24173.4]
  wire  tensorStore_io_vme_wr_data_ready; // @[Store.scala 52:27:@24173.4]
  wire  tensorStore_io_vme_wr_data_valid; // @[Store.scala 52:27:@24173.4]
  wire [63:0] tensorStore_io_vme_wr_data_bits; // @[Store.scala 52:27:@24173.4]
  wire  tensorStore_io_vme_wr_ack; // @[Store.scala 52:27:@24173.4]
  wire  tensorStore_io_tensor_wr_valid; // @[Store.scala 52:27:@24173.4]
  wire [10:0] tensorStore_io_tensor_wr_bits_idx; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_0; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_1; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_2; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_3; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_4; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_5; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_6; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_7; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_8; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_9; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_10; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_11; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_12; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_13; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_14; // @[Store.scala 52:27:@24173.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_15; // @[Store.scala 52:27:@24173.4]
  reg [1:0] state; // @[Store.scala 44:22:@24162.4]
  reg [31:0] _RAND_0;
  wire  _T_597; // @[Store.scala 54:40:@24176.4]
  wire  start; // @[Store.scala 54:35:@24177.4]
  wire  _T_598; // @[Conditional.scala 37:30:@24178.4]
  wire [1:0] _GEN_0; // @[Store.scala 63:36:@24185.10]
  wire [1:0] _GEN_1; // @[Store.scala 61:29:@24181.8]
  wire [1:0] _GEN_2; // @[Store.scala 60:19:@24180.6]
  wire  _T_599; // @[Conditional.scala 37:30:@24191.6]
  wire  _T_600; // @[Conditional.scala 37:30:@24196.8]
  wire [1:0] _GEN_3; // @[Store.scala 72:18:@24198.10]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@24197.8]
  wire [1:0] _GEN_5; // @[Conditional.scala 39:67:@24192.6]
  wire [1:0] _GEN_6; // @[Conditional.scala 40:58:@24179.4]
  wire  _T_601; // @[Store.scala 80:33:@24205.4]
  wire  _T_602; // @[Store.scala 80:42:@24206.4]
  wire  _T_603; // @[Store.scala 80:59:@24207.4]
  wire  _T_604; // @[Store.scala 80:50:@24208.4]
  wire  _T_605; // @[Store.scala 83:33:@24210.4]
  wire  _T_606; // @[Store.scala 83:43:@24211.4]
  Semaphore s ( // @[Store.scala 46:17:@24163.4]
    .clock(s_clock),
    .reset(s_reset),
    .io_spost(s_io_spost),
    .io_swait(s_io_swait),
    .io_sready(s_io_sready)
  );
  Queue_1 inst_q ( // @[Store.scala 47:22:@24166.4]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits)
  );
  StoreDecode dec ( // @[Store.scala 49:19:@24169.4]
    .io_inst(dec_io_inst),
    .io_push_prev(dec_io_push_prev),
    .io_pop_prev(dec_io_pop_prev),
    .io_isStore(dec_io_isStore),
    .io_isSync(dec_io_isSync)
  );
  TensorStore tensorStore ( // @[Store.scala 52:27:@24173.4]
    .clock(tensorStore_clock),
    .reset(tensorStore_reset),
    .io_start(tensorStore_io_start),
    .io_done(tensorStore_io_done),
    .io_inst(tensorStore_io_inst),
    .io_baddr(tensorStore_io_baddr),
    .io_vme_wr_cmd_ready(tensorStore_io_vme_wr_cmd_ready),
    .io_vme_wr_cmd_valid(tensorStore_io_vme_wr_cmd_valid),
    .io_vme_wr_cmd_bits_addr(tensorStore_io_vme_wr_cmd_bits_addr),
    .io_vme_wr_cmd_bits_len(tensorStore_io_vme_wr_cmd_bits_len),
    .io_vme_wr_data_ready(tensorStore_io_vme_wr_data_ready),
    .io_vme_wr_data_valid(tensorStore_io_vme_wr_data_valid),
    .io_vme_wr_data_bits(tensorStore_io_vme_wr_data_bits),
    .io_vme_wr_ack(tensorStore_io_vme_wr_ack),
    .io_tensor_wr_valid(tensorStore_io_tensor_wr_valid),
    .io_tensor_wr_bits_idx(tensorStore_io_tensor_wr_bits_idx),
    .io_tensor_wr_bits_data_0_0(tensorStore_io_tensor_wr_bits_data_0_0),
    .io_tensor_wr_bits_data_0_1(tensorStore_io_tensor_wr_bits_data_0_1),
    .io_tensor_wr_bits_data_0_2(tensorStore_io_tensor_wr_bits_data_0_2),
    .io_tensor_wr_bits_data_0_3(tensorStore_io_tensor_wr_bits_data_0_3),
    .io_tensor_wr_bits_data_0_4(tensorStore_io_tensor_wr_bits_data_0_4),
    .io_tensor_wr_bits_data_0_5(tensorStore_io_tensor_wr_bits_data_0_5),
    .io_tensor_wr_bits_data_0_6(tensorStore_io_tensor_wr_bits_data_0_6),
    .io_tensor_wr_bits_data_0_7(tensorStore_io_tensor_wr_bits_data_0_7),
    .io_tensor_wr_bits_data_0_8(tensorStore_io_tensor_wr_bits_data_0_8),
    .io_tensor_wr_bits_data_0_9(tensorStore_io_tensor_wr_bits_data_0_9),
    .io_tensor_wr_bits_data_0_10(tensorStore_io_tensor_wr_bits_data_0_10),
    .io_tensor_wr_bits_data_0_11(tensorStore_io_tensor_wr_bits_data_0_11),
    .io_tensor_wr_bits_data_0_12(tensorStore_io_tensor_wr_bits_data_0_12),
    .io_tensor_wr_bits_data_0_13(tensorStore_io_tensor_wr_bits_data_0_13),
    .io_tensor_wr_bits_data_0_14(tensorStore_io_tensor_wr_bits_data_0_14),
    .io_tensor_wr_bits_data_0_15(tensorStore_io_tensor_wr_bits_data_0_15)
  );
  assign _T_597 = dec_io_pop_prev ? s_io_sready : 1'h1; // @[Store.scala 54:40:@24176.4]
  assign start = inst_q_io_deq_valid & _T_597; // @[Store.scala 54:35:@24177.4]
  assign _T_598 = 2'h0 == state; // @[Conditional.scala 37:30:@24178.4]
  assign _GEN_0 = dec_io_isStore ? 2'h2 : state; // @[Store.scala 63:36:@24185.10]
  assign _GEN_1 = dec_io_isSync ? 2'h1 : _GEN_0; // @[Store.scala 61:29:@24181.8]
  assign _GEN_2 = start ? _GEN_1 : state; // @[Store.scala 60:19:@24180.6]
  assign _T_599 = 2'h1 == state; // @[Conditional.scala 37:30:@24191.6]
  assign _T_600 = 2'h2 == state; // @[Conditional.scala 37:30:@24196.8]
  assign _GEN_3 = tensorStore_io_done ? 2'h0 : state; // @[Store.scala 72:18:@24198.10]
  assign _GEN_4 = _T_600 ? _GEN_3 : state; // @[Conditional.scala 39:67:@24197.8]
  assign _GEN_5 = _T_599 ? 2'h0 : _GEN_4; // @[Conditional.scala 39:67:@24192.6]
  assign _GEN_6 = _T_598 ? _GEN_2 : _GEN_5; // @[Conditional.scala 40:58:@24179.4]
  assign _T_601 = state == 2'h2; // @[Store.scala 80:33:@24205.4]
  assign _T_602 = _T_601 & tensorStore_io_done; // @[Store.scala 80:42:@24206.4]
  assign _T_603 = state == 2'h1; // @[Store.scala 80:59:@24207.4]
  assign _T_604 = _T_602 | _T_603; // @[Store.scala 80:50:@24208.4]
  assign _T_605 = state == 2'h0; // @[Store.scala 83:33:@24210.4]
  assign _T_606 = _T_605 & start; // @[Store.scala 83:43:@24211.4]
  assign io_o_post = dec_io_push_prev & _T_604; // @[Store.scala 92:13:@24271.4]
  assign io_inst_ready = inst_q_io_enq_ready; // @[Store.scala 79:17:@24204.4]
  assign io_vme_wr_cmd_valid = tensorStore_io_vme_wr_cmd_valid; // @[Store.scala 86:13:@24222.4]
  assign io_vme_wr_cmd_bits_addr = tensorStore_io_vme_wr_cmd_bits_addr; // @[Store.scala 86:13:@24221.4]
  assign io_vme_wr_cmd_bits_len = tensorStore_io_vme_wr_cmd_bits_len; // @[Store.scala 86:13:@24220.4]
  assign io_vme_wr_data_valid = tensorStore_io_vme_wr_data_valid; // @[Store.scala 86:13:@24218.4]
  assign io_vme_wr_data_bits = tensorStore_io_vme_wr_data_bits; // @[Store.scala 86:13:@24217.4]
  assign s_clock = clock; // @[:@24164.4]
  assign s_reset = reset; // @[:@24165.4]
  assign s_io_spost = io_i_post; // @[Store.scala 90:14:@24261.4]
  assign s_io_swait = dec_io_pop_prev & _T_606; // @[Store.scala 91:14:@24265.4]
  assign inst_q_clock = clock; // @[:@24167.4]
  assign inst_q_reset = reset; // @[:@24168.4]
  assign inst_q_io_enq_valid = io_inst_valid; // @[Store.scala 79:17:@24203.4]
  assign inst_q_io_enq_bits = io_inst_bits; // @[Store.scala 79:17:@24202.4]
  assign inst_q_io_deq_ready = _T_602 | _T_603; // @[Store.scala 80:23:@24209.4]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Store.scala 50:15:@24172.4]
  assign tensorStore_clock = clock; // @[:@24174.4]
  assign tensorStore_reset = reset; // @[:@24175.4]
  assign tensorStore_io_start = _T_606 & dec_io_isStore; // @[Store.scala 83:24:@24213.4]
  assign tensorStore_io_inst = inst_q_io_deq_bits; // @[Store.scala 84:23:@24214.4]
  assign tensorStore_io_baddr = io_out_baddr; // @[Store.scala 85:24:@24215.4]
  assign tensorStore_io_vme_wr_cmd_ready = io_vme_wr_cmd_ready; // @[Store.scala 86:13:@24223.4]
  assign tensorStore_io_vme_wr_data_ready = io_vme_wr_data_ready; // @[Store.scala 86:13:@24219.4]
  assign tensorStore_io_vme_wr_ack = io_vme_wr_ack; // @[Store.scala 86:13:@24216.4]
  assign tensorStore_io_tensor_wr_valid = io_out_wr_valid; // @[Store.scala 87:25:@24241.4]
  assign tensorStore_io_tensor_wr_bits_idx = io_out_wr_bits_idx; // @[Store.scala 87:25:@24240.4]
  assign tensorStore_io_tensor_wr_bits_data_0_0 = io_out_wr_bits_data_0_0; // @[Store.scala 87:25:@24224.4]
  assign tensorStore_io_tensor_wr_bits_data_0_1 = io_out_wr_bits_data_0_1; // @[Store.scala 87:25:@24225.4]
  assign tensorStore_io_tensor_wr_bits_data_0_2 = io_out_wr_bits_data_0_2; // @[Store.scala 87:25:@24226.4]
  assign tensorStore_io_tensor_wr_bits_data_0_3 = io_out_wr_bits_data_0_3; // @[Store.scala 87:25:@24227.4]
  assign tensorStore_io_tensor_wr_bits_data_0_4 = io_out_wr_bits_data_0_4; // @[Store.scala 87:25:@24228.4]
  assign tensorStore_io_tensor_wr_bits_data_0_5 = io_out_wr_bits_data_0_5; // @[Store.scala 87:25:@24229.4]
  assign tensorStore_io_tensor_wr_bits_data_0_6 = io_out_wr_bits_data_0_6; // @[Store.scala 87:25:@24230.4]
  assign tensorStore_io_tensor_wr_bits_data_0_7 = io_out_wr_bits_data_0_7; // @[Store.scala 87:25:@24231.4]
  assign tensorStore_io_tensor_wr_bits_data_0_8 = io_out_wr_bits_data_0_8; // @[Store.scala 87:25:@24232.4]
  assign tensorStore_io_tensor_wr_bits_data_0_9 = io_out_wr_bits_data_0_9; // @[Store.scala 87:25:@24233.4]
  assign tensorStore_io_tensor_wr_bits_data_0_10 = io_out_wr_bits_data_0_10; // @[Store.scala 87:25:@24234.4]
  assign tensorStore_io_tensor_wr_bits_data_0_11 = io_out_wr_bits_data_0_11; // @[Store.scala 87:25:@24235.4]
  assign tensorStore_io_tensor_wr_bits_data_0_12 = io_out_wr_bits_data_0_12; // @[Store.scala 87:25:@24236.4]
  assign tensorStore_io_tensor_wr_bits_data_0_13 = io_out_wr_bits_data_0_13; // @[Store.scala 87:25:@24237.4]
  assign tensorStore_io_tensor_wr_bits_data_0_14 = io_out_wr_bits_data_0_14; // @[Store.scala 87:25:@24238.4]
  assign tensorStore_io_tensor_wr_bits_data_0_15 = io_out_wr_bits_data_0_15; // @[Store.scala 87:25:@24239.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_598) begin
        if (start) begin
          if (dec_io_isSync) begin
            state <= 2'h1;
          end else begin
            if (dec_io_isStore) begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_599) begin
          state <= 2'h0;
        end else begin
          if (_T_600) begin
            if (tensorStore_io_done) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module EventCounters( // @[:@24273.2]
  input         clock, // @[:@24274.4]
  input         reset, // @[:@24275.4]
  input         io_launch, // @[:@24276.4]
  input         io_finish, // @[:@24276.4]
  output        io_ecnt_0_valid, // @[:@24276.4]
  output [31:0] io_ecnt_0_bits, // @[:@24276.4]
  output        io_ucnt_0_valid, // @[:@24276.4]
  output [31:0] io_ucnt_0_bits, // @[:@24276.4]
  input         io_acc_wr_event // @[:@24276.4]
);
  reg [31:0] cycle_cnt; // @[EventCounters.scala 50:26:@24278.4]
  reg [31:0] _RAND_0;
  wire  _T_38; // @[EventCounters.scala 51:21:@24279.4]
  wire  _T_39; // @[EventCounters.scala 51:18:@24280.4]
  wire [32:0] _T_41; // @[EventCounters.scala 52:28:@24282.6]
  wire [31:0] _T_42; // @[EventCounters.scala 52:28:@24283.6]
  wire [31:0] _GEN_0; // @[EventCounters.scala 51:33:@24281.4]
  reg [31:0] acc_wr_count; // @[EventCounters.scala 59:25:@24291.4]
  reg [31:0] _RAND_1;
  wire  _T_46; // @[EventCounters.scala 60:9:@24292.4]
  wire  _T_47; // @[EventCounters.scala 60:20:@24293.4]
  wire [32:0] _T_50; // @[EventCounters.scala 63:34:@24299.8]
  wire [31:0] _T_51; // @[EventCounters.scala 63:34:@24300.8]
  wire [31:0] _GEN_1; // @[EventCounters.scala 62:32:@24298.6]
  assign _T_38 = io_finish == 1'h0; // @[EventCounters.scala 51:21:@24279.4]
  assign _T_39 = io_launch & _T_38; // @[EventCounters.scala 51:18:@24280.4]
  assign _T_41 = cycle_cnt + 32'h1; // @[EventCounters.scala 52:28:@24282.6]
  assign _T_42 = cycle_cnt + 32'h1; // @[EventCounters.scala 52:28:@24283.6]
  assign _GEN_0 = _T_39 ? _T_42 : 32'h0; // @[EventCounters.scala 51:33:@24281.4]
  assign _T_46 = io_launch == 1'h0; // @[EventCounters.scala 60:9:@24292.4]
  assign _T_47 = _T_46 | io_finish; // @[EventCounters.scala 60:20:@24293.4]
  assign _T_50 = acc_wr_count + 32'h1; // @[EventCounters.scala 63:34:@24299.8]
  assign _T_51 = acc_wr_count + 32'h1; // @[EventCounters.scala 63:34:@24300.8]
  assign _GEN_1 = io_acc_wr_event ? _T_51 : acc_wr_count; // @[EventCounters.scala 62:32:@24298.6]
  assign io_ecnt_0_valid = io_finish; // @[EventCounters.scala 56:20:@24289.4]
  assign io_ecnt_0_bits = cycle_cnt; // @[EventCounters.scala 57:19:@24290.4]
  assign io_ucnt_0_valid = io_finish; // @[EventCounters.scala 65:20:@24303.4]
  assign io_ucnt_0_bits = acc_wr_count; // @[EventCounters.scala 66:19:@24304.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycle_cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  acc_wr_count = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cycle_cnt <= 32'h0;
    end else begin
      if (_T_39) begin
        cycle_cnt <= _T_42;
      end else begin
        cycle_cnt <= 32'h0;
      end
    end
    if (_T_47) begin
      acc_wr_count <= 32'h0;
    end else begin
      if (io_acc_wr_event) begin
        acc_wr_count <= _T_51;
      end
    end
  end
endmodule
module Core( // @[:@24306.2]
  input         clock, // @[:@24307.4]
  input         reset, // @[:@24308.4]
  input         io_vcr_launch, // @[:@24309.4]
  output        io_vcr_finish, // @[:@24309.4]
  output        io_vcr_ecnt_0_valid, // @[:@24309.4]
  output [31:0] io_vcr_ecnt_0_bits, // @[:@24309.4]
  input  [31:0] io_vcr_vals_0, // @[:@24309.4]
  input  [31:0] io_vcr_ptrs_0, // @[:@24309.4]
  input  [31:0] io_vcr_ptrs_1, // @[:@24309.4]
  input  [31:0] io_vcr_ptrs_2, // @[:@24309.4]
  input  [31:0] io_vcr_ptrs_3, // @[:@24309.4]
  input  [31:0] io_vcr_ptrs_4, // @[:@24309.4]
  input  [31:0] io_vcr_ptrs_5, // @[:@24309.4]
  output        io_vcr_ucnt_0_valid, // @[:@24309.4]
  output [31:0] io_vcr_ucnt_0_bits, // @[:@24309.4]
  input         io_vme_rd_0_cmd_ready, // @[:@24309.4]
  output        io_vme_rd_0_cmd_valid, // @[:@24309.4]
  output [31:0] io_vme_rd_0_cmd_bits_addr, // @[:@24309.4]
  output [7:0]  io_vme_rd_0_cmd_bits_len, // @[:@24309.4]
  output        io_vme_rd_0_data_ready, // @[:@24309.4]
  input         io_vme_rd_0_data_valid, // @[:@24309.4]
  input  [63:0] io_vme_rd_0_data_bits, // @[:@24309.4]
  input         io_vme_rd_1_cmd_ready, // @[:@24309.4]
  output        io_vme_rd_1_cmd_valid, // @[:@24309.4]
  output [31:0] io_vme_rd_1_cmd_bits_addr, // @[:@24309.4]
  output [7:0]  io_vme_rd_1_cmd_bits_len, // @[:@24309.4]
  output        io_vme_rd_1_data_ready, // @[:@24309.4]
  input         io_vme_rd_1_data_valid, // @[:@24309.4]
  input  [63:0] io_vme_rd_1_data_bits, // @[:@24309.4]
  input         io_vme_rd_2_cmd_ready, // @[:@24309.4]
  output        io_vme_rd_2_cmd_valid, // @[:@24309.4]
  output [31:0] io_vme_rd_2_cmd_bits_addr, // @[:@24309.4]
  output [7:0]  io_vme_rd_2_cmd_bits_len, // @[:@24309.4]
  output        io_vme_rd_2_data_ready, // @[:@24309.4]
  input         io_vme_rd_2_data_valid, // @[:@24309.4]
  input  [63:0] io_vme_rd_2_data_bits, // @[:@24309.4]
  input         io_vme_rd_3_cmd_ready, // @[:@24309.4]
  output        io_vme_rd_3_cmd_valid, // @[:@24309.4]
  output [31:0] io_vme_rd_3_cmd_bits_addr, // @[:@24309.4]
  output [7:0]  io_vme_rd_3_cmd_bits_len, // @[:@24309.4]
  output        io_vme_rd_3_data_ready, // @[:@24309.4]
  input         io_vme_rd_3_data_valid, // @[:@24309.4]
  input  [63:0] io_vme_rd_3_data_bits, // @[:@24309.4]
  input         io_vme_rd_4_cmd_ready, // @[:@24309.4]
  output        io_vme_rd_4_cmd_valid, // @[:@24309.4]
  output [31:0] io_vme_rd_4_cmd_bits_addr, // @[:@24309.4]
  output [7:0]  io_vme_rd_4_cmd_bits_len, // @[:@24309.4]
  output        io_vme_rd_4_data_ready, // @[:@24309.4]
  input         io_vme_rd_4_data_valid, // @[:@24309.4]
  input  [63:0] io_vme_rd_4_data_bits, // @[:@24309.4]
  input         io_vme_wr_0_cmd_ready, // @[:@24309.4]
  output        io_vme_wr_0_cmd_valid, // @[:@24309.4]
  output [31:0] io_vme_wr_0_cmd_bits_addr, // @[:@24309.4]
  output [7:0]  io_vme_wr_0_cmd_bits_len, // @[:@24309.4]
  input         io_vme_wr_0_data_ready, // @[:@24309.4]
  output        io_vme_wr_0_data_valid, // @[:@24309.4]
  output [63:0] io_vme_wr_0_data_bits, // @[:@24309.4]
  input         io_vme_wr_0_ack // @[:@24309.4]
);
  wire  fetch_clock; // @[Core.scala 66:21:@24311.4]
  wire  fetch_reset; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_launch; // @[Core.scala 66:21:@24311.4]
  wire [31:0] fetch_io_ins_baddr; // @[Core.scala 66:21:@24311.4]
  wire [31:0] fetch_io_ins_count; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_vme_rd_cmd_ready; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_vme_rd_cmd_valid; // @[Core.scala 66:21:@24311.4]
  wire [31:0] fetch_io_vme_rd_cmd_bits_addr; // @[Core.scala 66:21:@24311.4]
  wire [7:0] fetch_io_vme_rd_cmd_bits_len; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_vme_rd_data_ready; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_vme_rd_data_valid; // @[Core.scala 66:21:@24311.4]
  wire [63:0] fetch_io_vme_rd_data_bits; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_inst_ld_ready; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_inst_ld_valid; // @[Core.scala 66:21:@24311.4]
  wire [127:0] fetch_io_inst_ld_bits; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_inst_co_ready; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_inst_co_valid; // @[Core.scala 66:21:@24311.4]
  wire [127:0] fetch_io_inst_co_bits; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_inst_st_ready; // @[Core.scala 66:21:@24311.4]
  wire  fetch_io_inst_st_valid; // @[Core.scala 66:21:@24311.4]
  wire [127:0] fetch_io_inst_st_bits; // @[Core.scala 66:21:@24311.4]
  wire  load_clock; // @[Core.scala 67:20:@24314.4]
  wire  load_reset; // @[Core.scala 67:20:@24314.4]
  wire  load_io_i_post; // @[Core.scala 67:20:@24314.4]
  wire  load_io_o_post; // @[Core.scala 67:20:@24314.4]
  wire  load_io_inst_ready; // @[Core.scala 67:20:@24314.4]
  wire  load_io_inst_valid; // @[Core.scala 67:20:@24314.4]
  wire [127:0] load_io_inst_bits; // @[Core.scala 67:20:@24314.4]
  wire [31:0] load_io_inp_baddr; // @[Core.scala 67:20:@24314.4]
  wire [31:0] load_io_wgt_baddr; // @[Core.scala 67:20:@24314.4]
  wire  load_io_vme_rd_0_cmd_ready; // @[Core.scala 67:20:@24314.4]
  wire  load_io_vme_rd_0_cmd_valid; // @[Core.scala 67:20:@24314.4]
  wire [31:0] load_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_vme_rd_0_cmd_bits_len; // @[Core.scala 67:20:@24314.4]
  wire  load_io_vme_rd_0_data_ready; // @[Core.scala 67:20:@24314.4]
  wire  load_io_vme_rd_0_data_valid; // @[Core.scala 67:20:@24314.4]
  wire [63:0] load_io_vme_rd_0_data_bits; // @[Core.scala 67:20:@24314.4]
  wire  load_io_vme_rd_1_cmd_ready; // @[Core.scala 67:20:@24314.4]
  wire  load_io_vme_rd_1_cmd_valid; // @[Core.scala 67:20:@24314.4]
  wire [31:0] load_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_vme_rd_1_cmd_bits_len; // @[Core.scala 67:20:@24314.4]
  wire  load_io_vme_rd_1_data_ready; // @[Core.scala 67:20:@24314.4]
  wire  load_io_vme_rd_1_data_valid; // @[Core.scala 67:20:@24314.4]
  wire [63:0] load_io_vme_rd_1_data_bits; // @[Core.scala 67:20:@24314.4]
  wire  load_io_inp_rd_idx_valid; // @[Core.scala 67:20:@24314.4]
  wire [10:0] load_io_inp_rd_idx_bits; // @[Core.scala 67:20:@24314.4]
  wire  load_io_inp_rd_data_valid; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_inp_rd_data_bits_0_15; // @[Core.scala 67:20:@24314.4]
  wire  load_io_wgt_rd_idx_valid; // @[Core.scala 67:20:@24314.4]
  wire [9:0] load_io_wgt_rd_idx_bits; // @[Core.scala 67:20:@24314.4]
  wire  load_io_wgt_rd_data_valid; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_15; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_0; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_1; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_2; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_3; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_4; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_5; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_6; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_7; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_8; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_9; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_10; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_11; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_12; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_13; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_14; // @[Core.scala 67:20:@24314.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_15; // @[Core.scala 67:20:@24314.4]
  wire  compute_clock; // @[Core.scala 68:23:@24317.4]
  wire  compute_reset; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_i_post_0; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_i_post_1; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_o_post_0; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_o_post_1; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_inst_ready; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_inst_valid; // @[Core.scala 68:23:@24317.4]
  wire [127:0] compute_io_inst_bits; // @[Core.scala 68:23:@24317.4]
  wire [31:0] compute_io_uop_baddr; // @[Core.scala 68:23:@24317.4]
  wire [31:0] compute_io_acc_baddr; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_vme_rd_0_cmd_ready; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_vme_rd_0_cmd_valid; // @[Core.scala 68:23:@24317.4]
  wire [31:0] compute_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_vme_rd_0_cmd_bits_len; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_vme_rd_0_data_ready; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_vme_rd_0_data_valid; // @[Core.scala 68:23:@24317.4]
  wire [63:0] compute_io_vme_rd_0_data_bits; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_vme_rd_1_cmd_ready; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_vme_rd_1_cmd_valid; // @[Core.scala 68:23:@24317.4]
  wire [31:0] compute_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_vme_rd_1_cmd_bits_len; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_vme_rd_1_data_ready; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_vme_rd_1_data_valid; // @[Core.scala 68:23:@24317.4]
  wire [63:0] compute_io_vme_rd_1_data_bits; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_inp_rd_idx_valid; // @[Core.scala 68:23:@24317.4]
  wire [10:0] compute_io_inp_rd_idx_bits; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_inp_rd_data_valid; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_15; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_wgt_rd_idx_valid; // @[Core.scala 68:23:@24317.4]
  wire [9:0] compute_io_wgt_rd_idx_bits; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_wgt_rd_data_valid; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_15; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_15; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_out_wr_valid; // @[Core.scala 68:23:@24317.4]
  wire [10:0] compute_io_out_wr_bits_idx; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_0; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_1; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_2; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_3; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_4; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_5; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_6; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_7; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_8; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_9; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_10; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_11; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_12; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_13; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_14; // @[Core.scala 68:23:@24317.4]
  wire [7:0] compute_io_out_wr_bits_data_0_15; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_finish; // @[Core.scala 68:23:@24317.4]
  wire  compute_io_acc_wr_event; // @[Core.scala 68:23:@24317.4]
  wire  store_clock; // @[Core.scala 69:21:@24320.4]
  wire  store_reset; // @[Core.scala 69:21:@24320.4]
  wire  store_io_i_post; // @[Core.scala 69:21:@24320.4]
  wire  store_io_o_post; // @[Core.scala 69:21:@24320.4]
  wire  store_io_inst_ready; // @[Core.scala 69:21:@24320.4]
  wire  store_io_inst_valid; // @[Core.scala 69:21:@24320.4]
  wire [127:0] store_io_inst_bits; // @[Core.scala 69:21:@24320.4]
  wire [31:0] store_io_out_baddr; // @[Core.scala 69:21:@24320.4]
  wire  store_io_vme_wr_cmd_ready; // @[Core.scala 69:21:@24320.4]
  wire  store_io_vme_wr_cmd_valid; // @[Core.scala 69:21:@24320.4]
  wire [31:0] store_io_vme_wr_cmd_bits_addr; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_vme_wr_cmd_bits_len; // @[Core.scala 69:21:@24320.4]
  wire  store_io_vme_wr_data_ready; // @[Core.scala 69:21:@24320.4]
  wire  store_io_vme_wr_data_valid; // @[Core.scala 69:21:@24320.4]
  wire [63:0] store_io_vme_wr_data_bits; // @[Core.scala 69:21:@24320.4]
  wire  store_io_vme_wr_ack; // @[Core.scala 69:21:@24320.4]
  wire  store_io_out_wr_valid; // @[Core.scala 69:21:@24320.4]
  wire [10:0] store_io_out_wr_bits_idx; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_0; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_1; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_2; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_3; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_4; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_5; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_6; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_7; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_8; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_9; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_10; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_11; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_12; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_13; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_14; // @[Core.scala 69:21:@24320.4]
  wire [7:0] store_io_out_wr_bits_data_0_15; // @[Core.scala 69:21:@24320.4]
  wire  ecounters_clock; // @[Core.scala 70:25:@24323.4]
  wire  ecounters_reset; // @[Core.scala 70:25:@24323.4]
  wire  ecounters_io_launch; // @[Core.scala 70:25:@24323.4]
  wire  ecounters_io_finish; // @[Core.scala 70:25:@24323.4]
  wire  ecounters_io_ecnt_0_valid; // @[Core.scala 70:25:@24323.4]
  wire [31:0] ecounters_io_ecnt_0_bits; // @[Core.scala 70:25:@24323.4]
  wire  ecounters_io_ucnt_0_valid; // @[Core.scala 70:25:@24323.4]
  wire [31:0] ecounters_io_ucnt_0_bits; // @[Core.scala 70:25:@24323.4]
  wire  ecounters_io_acc_wr_event; // @[Core.scala 70:25:@24323.4]
  reg  finish; // @[Core.scala 118:23:@24988.4]
  reg [31:0] _RAND_0;
  Fetch fetch ( // @[Core.scala 66:21:@24311.4]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_launch(fetch_io_launch),
    .io_ins_baddr(fetch_io_ins_baddr),
    .io_ins_count(fetch_io_ins_count),
    .io_vme_rd_cmd_ready(fetch_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(fetch_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(fetch_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(fetch_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(fetch_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(fetch_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(fetch_io_vme_rd_data_bits),
    .io_inst_ld_ready(fetch_io_inst_ld_ready),
    .io_inst_ld_valid(fetch_io_inst_ld_valid),
    .io_inst_ld_bits(fetch_io_inst_ld_bits),
    .io_inst_co_ready(fetch_io_inst_co_ready),
    .io_inst_co_valid(fetch_io_inst_co_valid),
    .io_inst_co_bits(fetch_io_inst_co_bits),
    .io_inst_st_ready(fetch_io_inst_st_ready),
    .io_inst_st_valid(fetch_io_inst_st_valid),
    .io_inst_st_bits(fetch_io_inst_st_bits)
  );
  Load load ( // @[Core.scala 67:20:@24314.4]
    .clock(load_clock),
    .reset(load_reset),
    .io_i_post(load_io_i_post),
    .io_o_post(load_io_o_post),
    .io_inst_ready(load_io_inst_ready),
    .io_inst_valid(load_io_inst_valid),
    .io_inst_bits(load_io_inst_bits),
    .io_inp_baddr(load_io_inp_baddr),
    .io_wgt_baddr(load_io_wgt_baddr),
    .io_vme_rd_0_cmd_ready(load_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(load_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(load_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(load_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(load_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(load_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits(load_io_vme_rd_0_data_bits),
    .io_vme_rd_1_cmd_ready(load_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(load_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(load_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(load_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_data_ready(load_io_vme_rd_1_data_ready),
    .io_vme_rd_1_data_valid(load_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits(load_io_vme_rd_1_data_bits),
    .io_inp_rd_idx_valid(load_io_inp_rd_idx_valid),
    .io_inp_rd_idx_bits(load_io_inp_rd_idx_bits),
    .io_inp_rd_data_valid(load_io_inp_rd_data_valid),
    .io_inp_rd_data_bits_0_0(load_io_inp_rd_data_bits_0_0),
    .io_inp_rd_data_bits_0_1(load_io_inp_rd_data_bits_0_1),
    .io_inp_rd_data_bits_0_2(load_io_inp_rd_data_bits_0_2),
    .io_inp_rd_data_bits_0_3(load_io_inp_rd_data_bits_0_3),
    .io_inp_rd_data_bits_0_4(load_io_inp_rd_data_bits_0_4),
    .io_inp_rd_data_bits_0_5(load_io_inp_rd_data_bits_0_5),
    .io_inp_rd_data_bits_0_6(load_io_inp_rd_data_bits_0_6),
    .io_inp_rd_data_bits_0_7(load_io_inp_rd_data_bits_0_7),
    .io_inp_rd_data_bits_0_8(load_io_inp_rd_data_bits_0_8),
    .io_inp_rd_data_bits_0_9(load_io_inp_rd_data_bits_0_9),
    .io_inp_rd_data_bits_0_10(load_io_inp_rd_data_bits_0_10),
    .io_inp_rd_data_bits_0_11(load_io_inp_rd_data_bits_0_11),
    .io_inp_rd_data_bits_0_12(load_io_inp_rd_data_bits_0_12),
    .io_inp_rd_data_bits_0_13(load_io_inp_rd_data_bits_0_13),
    .io_inp_rd_data_bits_0_14(load_io_inp_rd_data_bits_0_14),
    .io_inp_rd_data_bits_0_15(load_io_inp_rd_data_bits_0_15),
    .io_wgt_rd_idx_valid(load_io_wgt_rd_idx_valid),
    .io_wgt_rd_idx_bits(load_io_wgt_rd_idx_bits),
    .io_wgt_rd_data_valid(load_io_wgt_rd_data_valid),
    .io_wgt_rd_data_bits_0_0(load_io_wgt_rd_data_bits_0_0),
    .io_wgt_rd_data_bits_0_1(load_io_wgt_rd_data_bits_0_1),
    .io_wgt_rd_data_bits_0_2(load_io_wgt_rd_data_bits_0_2),
    .io_wgt_rd_data_bits_0_3(load_io_wgt_rd_data_bits_0_3),
    .io_wgt_rd_data_bits_0_4(load_io_wgt_rd_data_bits_0_4),
    .io_wgt_rd_data_bits_0_5(load_io_wgt_rd_data_bits_0_5),
    .io_wgt_rd_data_bits_0_6(load_io_wgt_rd_data_bits_0_6),
    .io_wgt_rd_data_bits_0_7(load_io_wgt_rd_data_bits_0_7),
    .io_wgt_rd_data_bits_0_8(load_io_wgt_rd_data_bits_0_8),
    .io_wgt_rd_data_bits_0_9(load_io_wgt_rd_data_bits_0_9),
    .io_wgt_rd_data_bits_0_10(load_io_wgt_rd_data_bits_0_10),
    .io_wgt_rd_data_bits_0_11(load_io_wgt_rd_data_bits_0_11),
    .io_wgt_rd_data_bits_0_12(load_io_wgt_rd_data_bits_0_12),
    .io_wgt_rd_data_bits_0_13(load_io_wgt_rd_data_bits_0_13),
    .io_wgt_rd_data_bits_0_14(load_io_wgt_rd_data_bits_0_14),
    .io_wgt_rd_data_bits_0_15(load_io_wgt_rd_data_bits_0_15),
    .io_wgt_rd_data_bits_1_0(load_io_wgt_rd_data_bits_1_0),
    .io_wgt_rd_data_bits_1_1(load_io_wgt_rd_data_bits_1_1),
    .io_wgt_rd_data_bits_1_2(load_io_wgt_rd_data_bits_1_2),
    .io_wgt_rd_data_bits_1_3(load_io_wgt_rd_data_bits_1_3),
    .io_wgt_rd_data_bits_1_4(load_io_wgt_rd_data_bits_1_4),
    .io_wgt_rd_data_bits_1_5(load_io_wgt_rd_data_bits_1_5),
    .io_wgt_rd_data_bits_1_6(load_io_wgt_rd_data_bits_1_6),
    .io_wgt_rd_data_bits_1_7(load_io_wgt_rd_data_bits_1_7),
    .io_wgt_rd_data_bits_1_8(load_io_wgt_rd_data_bits_1_8),
    .io_wgt_rd_data_bits_1_9(load_io_wgt_rd_data_bits_1_9),
    .io_wgt_rd_data_bits_1_10(load_io_wgt_rd_data_bits_1_10),
    .io_wgt_rd_data_bits_1_11(load_io_wgt_rd_data_bits_1_11),
    .io_wgt_rd_data_bits_1_12(load_io_wgt_rd_data_bits_1_12),
    .io_wgt_rd_data_bits_1_13(load_io_wgt_rd_data_bits_1_13),
    .io_wgt_rd_data_bits_1_14(load_io_wgt_rd_data_bits_1_14),
    .io_wgt_rd_data_bits_1_15(load_io_wgt_rd_data_bits_1_15),
    .io_wgt_rd_data_bits_2_0(load_io_wgt_rd_data_bits_2_0),
    .io_wgt_rd_data_bits_2_1(load_io_wgt_rd_data_bits_2_1),
    .io_wgt_rd_data_bits_2_2(load_io_wgt_rd_data_bits_2_2),
    .io_wgt_rd_data_bits_2_3(load_io_wgt_rd_data_bits_2_3),
    .io_wgt_rd_data_bits_2_4(load_io_wgt_rd_data_bits_2_4),
    .io_wgt_rd_data_bits_2_5(load_io_wgt_rd_data_bits_2_5),
    .io_wgt_rd_data_bits_2_6(load_io_wgt_rd_data_bits_2_6),
    .io_wgt_rd_data_bits_2_7(load_io_wgt_rd_data_bits_2_7),
    .io_wgt_rd_data_bits_2_8(load_io_wgt_rd_data_bits_2_8),
    .io_wgt_rd_data_bits_2_9(load_io_wgt_rd_data_bits_2_9),
    .io_wgt_rd_data_bits_2_10(load_io_wgt_rd_data_bits_2_10),
    .io_wgt_rd_data_bits_2_11(load_io_wgt_rd_data_bits_2_11),
    .io_wgt_rd_data_bits_2_12(load_io_wgt_rd_data_bits_2_12),
    .io_wgt_rd_data_bits_2_13(load_io_wgt_rd_data_bits_2_13),
    .io_wgt_rd_data_bits_2_14(load_io_wgt_rd_data_bits_2_14),
    .io_wgt_rd_data_bits_2_15(load_io_wgt_rd_data_bits_2_15),
    .io_wgt_rd_data_bits_3_0(load_io_wgt_rd_data_bits_3_0),
    .io_wgt_rd_data_bits_3_1(load_io_wgt_rd_data_bits_3_1),
    .io_wgt_rd_data_bits_3_2(load_io_wgt_rd_data_bits_3_2),
    .io_wgt_rd_data_bits_3_3(load_io_wgt_rd_data_bits_3_3),
    .io_wgt_rd_data_bits_3_4(load_io_wgt_rd_data_bits_3_4),
    .io_wgt_rd_data_bits_3_5(load_io_wgt_rd_data_bits_3_5),
    .io_wgt_rd_data_bits_3_6(load_io_wgt_rd_data_bits_3_6),
    .io_wgt_rd_data_bits_3_7(load_io_wgt_rd_data_bits_3_7),
    .io_wgt_rd_data_bits_3_8(load_io_wgt_rd_data_bits_3_8),
    .io_wgt_rd_data_bits_3_9(load_io_wgt_rd_data_bits_3_9),
    .io_wgt_rd_data_bits_3_10(load_io_wgt_rd_data_bits_3_10),
    .io_wgt_rd_data_bits_3_11(load_io_wgt_rd_data_bits_3_11),
    .io_wgt_rd_data_bits_3_12(load_io_wgt_rd_data_bits_3_12),
    .io_wgt_rd_data_bits_3_13(load_io_wgt_rd_data_bits_3_13),
    .io_wgt_rd_data_bits_3_14(load_io_wgt_rd_data_bits_3_14),
    .io_wgt_rd_data_bits_3_15(load_io_wgt_rd_data_bits_3_15),
    .io_wgt_rd_data_bits_4_0(load_io_wgt_rd_data_bits_4_0),
    .io_wgt_rd_data_bits_4_1(load_io_wgt_rd_data_bits_4_1),
    .io_wgt_rd_data_bits_4_2(load_io_wgt_rd_data_bits_4_2),
    .io_wgt_rd_data_bits_4_3(load_io_wgt_rd_data_bits_4_3),
    .io_wgt_rd_data_bits_4_4(load_io_wgt_rd_data_bits_4_4),
    .io_wgt_rd_data_bits_4_5(load_io_wgt_rd_data_bits_4_5),
    .io_wgt_rd_data_bits_4_6(load_io_wgt_rd_data_bits_4_6),
    .io_wgt_rd_data_bits_4_7(load_io_wgt_rd_data_bits_4_7),
    .io_wgt_rd_data_bits_4_8(load_io_wgt_rd_data_bits_4_8),
    .io_wgt_rd_data_bits_4_9(load_io_wgt_rd_data_bits_4_9),
    .io_wgt_rd_data_bits_4_10(load_io_wgt_rd_data_bits_4_10),
    .io_wgt_rd_data_bits_4_11(load_io_wgt_rd_data_bits_4_11),
    .io_wgt_rd_data_bits_4_12(load_io_wgt_rd_data_bits_4_12),
    .io_wgt_rd_data_bits_4_13(load_io_wgt_rd_data_bits_4_13),
    .io_wgt_rd_data_bits_4_14(load_io_wgt_rd_data_bits_4_14),
    .io_wgt_rd_data_bits_4_15(load_io_wgt_rd_data_bits_4_15),
    .io_wgt_rd_data_bits_5_0(load_io_wgt_rd_data_bits_5_0),
    .io_wgt_rd_data_bits_5_1(load_io_wgt_rd_data_bits_5_1),
    .io_wgt_rd_data_bits_5_2(load_io_wgt_rd_data_bits_5_2),
    .io_wgt_rd_data_bits_5_3(load_io_wgt_rd_data_bits_5_3),
    .io_wgt_rd_data_bits_5_4(load_io_wgt_rd_data_bits_5_4),
    .io_wgt_rd_data_bits_5_5(load_io_wgt_rd_data_bits_5_5),
    .io_wgt_rd_data_bits_5_6(load_io_wgt_rd_data_bits_5_6),
    .io_wgt_rd_data_bits_5_7(load_io_wgt_rd_data_bits_5_7),
    .io_wgt_rd_data_bits_5_8(load_io_wgt_rd_data_bits_5_8),
    .io_wgt_rd_data_bits_5_9(load_io_wgt_rd_data_bits_5_9),
    .io_wgt_rd_data_bits_5_10(load_io_wgt_rd_data_bits_5_10),
    .io_wgt_rd_data_bits_5_11(load_io_wgt_rd_data_bits_5_11),
    .io_wgt_rd_data_bits_5_12(load_io_wgt_rd_data_bits_5_12),
    .io_wgt_rd_data_bits_5_13(load_io_wgt_rd_data_bits_5_13),
    .io_wgt_rd_data_bits_5_14(load_io_wgt_rd_data_bits_5_14),
    .io_wgt_rd_data_bits_5_15(load_io_wgt_rd_data_bits_5_15),
    .io_wgt_rd_data_bits_6_0(load_io_wgt_rd_data_bits_6_0),
    .io_wgt_rd_data_bits_6_1(load_io_wgt_rd_data_bits_6_1),
    .io_wgt_rd_data_bits_6_2(load_io_wgt_rd_data_bits_6_2),
    .io_wgt_rd_data_bits_6_3(load_io_wgt_rd_data_bits_6_3),
    .io_wgt_rd_data_bits_6_4(load_io_wgt_rd_data_bits_6_4),
    .io_wgt_rd_data_bits_6_5(load_io_wgt_rd_data_bits_6_5),
    .io_wgt_rd_data_bits_6_6(load_io_wgt_rd_data_bits_6_6),
    .io_wgt_rd_data_bits_6_7(load_io_wgt_rd_data_bits_6_7),
    .io_wgt_rd_data_bits_6_8(load_io_wgt_rd_data_bits_6_8),
    .io_wgt_rd_data_bits_6_9(load_io_wgt_rd_data_bits_6_9),
    .io_wgt_rd_data_bits_6_10(load_io_wgt_rd_data_bits_6_10),
    .io_wgt_rd_data_bits_6_11(load_io_wgt_rd_data_bits_6_11),
    .io_wgt_rd_data_bits_6_12(load_io_wgt_rd_data_bits_6_12),
    .io_wgt_rd_data_bits_6_13(load_io_wgt_rd_data_bits_6_13),
    .io_wgt_rd_data_bits_6_14(load_io_wgt_rd_data_bits_6_14),
    .io_wgt_rd_data_bits_6_15(load_io_wgt_rd_data_bits_6_15),
    .io_wgt_rd_data_bits_7_0(load_io_wgt_rd_data_bits_7_0),
    .io_wgt_rd_data_bits_7_1(load_io_wgt_rd_data_bits_7_1),
    .io_wgt_rd_data_bits_7_2(load_io_wgt_rd_data_bits_7_2),
    .io_wgt_rd_data_bits_7_3(load_io_wgt_rd_data_bits_7_3),
    .io_wgt_rd_data_bits_7_4(load_io_wgt_rd_data_bits_7_4),
    .io_wgt_rd_data_bits_7_5(load_io_wgt_rd_data_bits_7_5),
    .io_wgt_rd_data_bits_7_6(load_io_wgt_rd_data_bits_7_6),
    .io_wgt_rd_data_bits_7_7(load_io_wgt_rd_data_bits_7_7),
    .io_wgt_rd_data_bits_7_8(load_io_wgt_rd_data_bits_7_8),
    .io_wgt_rd_data_bits_7_9(load_io_wgt_rd_data_bits_7_9),
    .io_wgt_rd_data_bits_7_10(load_io_wgt_rd_data_bits_7_10),
    .io_wgt_rd_data_bits_7_11(load_io_wgt_rd_data_bits_7_11),
    .io_wgt_rd_data_bits_7_12(load_io_wgt_rd_data_bits_7_12),
    .io_wgt_rd_data_bits_7_13(load_io_wgt_rd_data_bits_7_13),
    .io_wgt_rd_data_bits_7_14(load_io_wgt_rd_data_bits_7_14),
    .io_wgt_rd_data_bits_7_15(load_io_wgt_rd_data_bits_7_15),
    .io_wgt_rd_data_bits_8_0(load_io_wgt_rd_data_bits_8_0),
    .io_wgt_rd_data_bits_8_1(load_io_wgt_rd_data_bits_8_1),
    .io_wgt_rd_data_bits_8_2(load_io_wgt_rd_data_bits_8_2),
    .io_wgt_rd_data_bits_8_3(load_io_wgt_rd_data_bits_8_3),
    .io_wgt_rd_data_bits_8_4(load_io_wgt_rd_data_bits_8_4),
    .io_wgt_rd_data_bits_8_5(load_io_wgt_rd_data_bits_8_5),
    .io_wgt_rd_data_bits_8_6(load_io_wgt_rd_data_bits_8_6),
    .io_wgt_rd_data_bits_8_7(load_io_wgt_rd_data_bits_8_7),
    .io_wgt_rd_data_bits_8_8(load_io_wgt_rd_data_bits_8_8),
    .io_wgt_rd_data_bits_8_9(load_io_wgt_rd_data_bits_8_9),
    .io_wgt_rd_data_bits_8_10(load_io_wgt_rd_data_bits_8_10),
    .io_wgt_rd_data_bits_8_11(load_io_wgt_rd_data_bits_8_11),
    .io_wgt_rd_data_bits_8_12(load_io_wgt_rd_data_bits_8_12),
    .io_wgt_rd_data_bits_8_13(load_io_wgt_rd_data_bits_8_13),
    .io_wgt_rd_data_bits_8_14(load_io_wgt_rd_data_bits_8_14),
    .io_wgt_rd_data_bits_8_15(load_io_wgt_rd_data_bits_8_15),
    .io_wgt_rd_data_bits_9_0(load_io_wgt_rd_data_bits_9_0),
    .io_wgt_rd_data_bits_9_1(load_io_wgt_rd_data_bits_9_1),
    .io_wgt_rd_data_bits_9_2(load_io_wgt_rd_data_bits_9_2),
    .io_wgt_rd_data_bits_9_3(load_io_wgt_rd_data_bits_9_3),
    .io_wgt_rd_data_bits_9_4(load_io_wgt_rd_data_bits_9_4),
    .io_wgt_rd_data_bits_9_5(load_io_wgt_rd_data_bits_9_5),
    .io_wgt_rd_data_bits_9_6(load_io_wgt_rd_data_bits_9_6),
    .io_wgt_rd_data_bits_9_7(load_io_wgt_rd_data_bits_9_7),
    .io_wgt_rd_data_bits_9_8(load_io_wgt_rd_data_bits_9_8),
    .io_wgt_rd_data_bits_9_9(load_io_wgt_rd_data_bits_9_9),
    .io_wgt_rd_data_bits_9_10(load_io_wgt_rd_data_bits_9_10),
    .io_wgt_rd_data_bits_9_11(load_io_wgt_rd_data_bits_9_11),
    .io_wgt_rd_data_bits_9_12(load_io_wgt_rd_data_bits_9_12),
    .io_wgt_rd_data_bits_9_13(load_io_wgt_rd_data_bits_9_13),
    .io_wgt_rd_data_bits_9_14(load_io_wgt_rd_data_bits_9_14),
    .io_wgt_rd_data_bits_9_15(load_io_wgt_rd_data_bits_9_15),
    .io_wgt_rd_data_bits_10_0(load_io_wgt_rd_data_bits_10_0),
    .io_wgt_rd_data_bits_10_1(load_io_wgt_rd_data_bits_10_1),
    .io_wgt_rd_data_bits_10_2(load_io_wgt_rd_data_bits_10_2),
    .io_wgt_rd_data_bits_10_3(load_io_wgt_rd_data_bits_10_3),
    .io_wgt_rd_data_bits_10_4(load_io_wgt_rd_data_bits_10_4),
    .io_wgt_rd_data_bits_10_5(load_io_wgt_rd_data_bits_10_5),
    .io_wgt_rd_data_bits_10_6(load_io_wgt_rd_data_bits_10_6),
    .io_wgt_rd_data_bits_10_7(load_io_wgt_rd_data_bits_10_7),
    .io_wgt_rd_data_bits_10_8(load_io_wgt_rd_data_bits_10_8),
    .io_wgt_rd_data_bits_10_9(load_io_wgt_rd_data_bits_10_9),
    .io_wgt_rd_data_bits_10_10(load_io_wgt_rd_data_bits_10_10),
    .io_wgt_rd_data_bits_10_11(load_io_wgt_rd_data_bits_10_11),
    .io_wgt_rd_data_bits_10_12(load_io_wgt_rd_data_bits_10_12),
    .io_wgt_rd_data_bits_10_13(load_io_wgt_rd_data_bits_10_13),
    .io_wgt_rd_data_bits_10_14(load_io_wgt_rd_data_bits_10_14),
    .io_wgt_rd_data_bits_10_15(load_io_wgt_rd_data_bits_10_15),
    .io_wgt_rd_data_bits_11_0(load_io_wgt_rd_data_bits_11_0),
    .io_wgt_rd_data_bits_11_1(load_io_wgt_rd_data_bits_11_1),
    .io_wgt_rd_data_bits_11_2(load_io_wgt_rd_data_bits_11_2),
    .io_wgt_rd_data_bits_11_3(load_io_wgt_rd_data_bits_11_3),
    .io_wgt_rd_data_bits_11_4(load_io_wgt_rd_data_bits_11_4),
    .io_wgt_rd_data_bits_11_5(load_io_wgt_rd_data_bits_11_5),
    .io_wgt_rd_data_bits_11_6(load_io_wgt_rd_data_bits_11_6),
    .io_wgt_rd_data_bits_11_7(load_io_wgt_rd_data_bits_11_7),
    .io_wgt_rd_data_bits_11_8(load_io_wgt_rd_data_bits_11_8),
    .io_wgt_rd_data_bits_11_9(load_io_wgt_rd_data_bits_11_9),
    .io_wgt_rd_data_bits_11_10(load_io_wgt_rd_data_bits_11_10),
    .io_wgt_rd_data_bits_11_11(load_io_wgt_rd_data_bits_11_11),
    .io_wgt_rd_data_bits_11_12(load_io_wgt_rd_data_bits_11_12),
    .io_wgt_rd_data_bits_11_13(load_io_wgt_rd_data_bits_11_13),
    .io_wgt_rd_data_bits_11_14(load_io_wgt_rd_data_bits_11_14),
    .io_wgt_rd_data_bits_11_15(load_io_wgt_rd_data_bits_11_15),
    .io_wgt_rd_data_bits_12_0(load_io_wgt_rd_data_bits_12_0),
    .io_wgt_rd_data_bits_12_1(load_io_wgt_rd_data_bits_12_1),
    .io_wgt_rd_data_bits_12_2(load_io_wgt_rd_data_bits_12_2),
    .io_wgt_rd_data_bits_12_3(load_io_wgt_rd_data_bits_12_3),
    .io_wgt_rd_data_bits_12_4(load_io_wgt_rd_data_bits_12_4),
    .io_wgt_rd_data_bits_12_5(load_io_wgt_rd_data_bits_12_5),
    .io_wgt_rd_data_bits_12_6(load_io_wgt_rd_data_bits_12_6),
    .io_wgt_rd_data_bits_12_7(load_io_wgt_rd_data_bits_12_7),
    .io_wgt_rd_data_bits_12_8(load_io_wgt_rd_data_bits_12_8),
    .io_wgt_rd_data_bits_12_9(load_io_wgt_rd_data_bits_12_9),
    .io_wgt_rd_data_bits_12_10(load_io_wgt_rd_data_bits_12_10),
    .io_wgt_rd_data_bits_12_11(load_io_wgt_rd_data_bits_12_11),
    .io_wgt_rd_data_bits_12_12(load_io_wgt_rd_data_bits_12_12),
    .io_wgt_rd_data_bits_12_13(load_io_wgt_rd_data_bits_12_13),
    .io_wgt_rd_data_bits_12_14(load_io_wgt_rd_data_bits_12_14),
    .io_wgt_rd_data_bits_12_15(load_io_wgt_rd_data_bits_12_15),
    .io_wgt_rd_data_bits_13_0(load_io_wgt_rd_data_bits_13_0),
    .io_wgt_rd_data_bits_13_1(load_io_wgt_rd_data_bits_13_1),
    .io_wgt_rd_data_bits_13_2(load_io_wgt_rd_data_bits_13_2),
    .io_wgt_rd_data_bits_13_3(load_io_wgt_rd_data_bits_13_3),
    .io_wgt_rd_data_bits_13_4(load_io_wgt_rd_data_bits_13_4),
    .io_wgt_rd_data_bits_13_5(load_io_wgt_rd_data_bits_13_5),
    .io_wgt_rd_data_bits_13_6(load_io_wgt_rd_data_bits_13_6),
    .io_wgt_rd_data_bits_13_7(load_io_wgt_rd_data_bits_13_7),
    .io_wgt_rd_data_bits_13_8(load_io_wgt_rd_data_bits_13_8),
    .io_wgt_rd_data_bits_13_9(load_io_wgt_rd_data_bits_13_9),
    .io_wgt_rd_data_bits_13_10(load_io_wgt_rd_data_bits_13_10),
    .io_wgt_rd_data_bits_13_11(load_io_wgt_rd_data_bits_13_11),
    .io_wgt_rd_data_bits_13_12(load_io_wgt_rd_data_bits_13_12),
    .io_wgt_rd_data_bits_13_13(load_io_wgt_rd_data_bits_13_13),
    .io_wgt_rd_data_bits_13_14(load_io_wgt_rd_data_bits_13_14),
    .io_wgt_rd_data_bits_13_15(load_io_wgt_rd_data_bits_13_15),
    .io_wgt_rd_data_bits_14_0(load_io_wgt_rd_data_bits_14_0),
    .io_wgt_rd_data_bits_14_1(load_io_wgt_rd_data_bits_14_1),
    .io_wgt_rd_data_bits_14_2(load_io_wgt_rd_data_bits_14_2),
    .io_wgt_rd_data_bits_14_3(load_io_wgt_rd_data_bits_14_3),
    .io_wgt_rd_data_bits_14_4(load_io_wgt_rd_data_bits_14_4),
    .io_wgt_rd_data_bits_14_5(load_io_wgt_rd_data_bits_14_5),
    .io_wgt_rd_data_bits_14_6(load_io_wgt_rd_data_bits_14_6),
    .io_wgt_rd_data_bits_14_7(load_io_wgt_rd_data_bits_14_7),
    .io_wgt_rd_data_bits_14_8(load_io_wgt_rd_data_bits_14_8),
    .io_wgt_rd_data_bits_14_9(load_io_wgt_rd_data_bits_14_9),
    .io_wgt_rd_data_bits_14_10(load_io_wgt_rd_data_bits_14_10),
    .io_wgt_rd_data_bits_14_11(load_io_wgt_rd_data_bits_14_11),
    .io_wgt_rd_data_bits_14_12(load_io_wgt_rd_data_bits_14_12),
    .io_wgt_rd_data_bits_14_13(load_io_wgt_rd_data_bits_14_13),
    .io_wgt_rd_data_bits_14_14(load_io_wgt_rd_data_bits_14_14),
    .io_wgt_rd_data_bits_14_15(load_io_wgt_rd_data_bits_14_15),
    .io_wgt_rd_data_bits_15_0(load_io_wgt_rd_data_bits_15_0),
    .io_wgt_rd_data_bits_15_1(load_io_wgt_rd_data_bits_15_1),
    .io_wgt_rd_data_bits_15_2(load_io_wgt_rd_data_bits_15_2),
    .io_wgt_rd_data_bits_15_3(load_io_wgt_rd_data_bits_15_3),
    .io_wgt_rd_data_bits_15_4(load_io_wgt_rd_data_bits_15_4),
    .io_wgt_rd_data_bits_15_5(load_io_wgt_rd_data_bits_15_5),
    .io_wgt_rd_data_bits_15_6(load_io_wgt_rd_data_bits_15_6),
    .io_wgt_rd_data_bits_15_7(load_io_wgt_rd_data_bits_15_7),
    .io_wgt_rd_data_bits_15_8(load_io_wgt_rd_data_bits_15_8),
    .io_wgt_rd_data_bits_15_9(load_io_wgt_rd_data_bits_15_9),
    .io_wgt_rd_data_bits_15_10(load_io_wgt_rd_data_bits_15_10),
    .io_wgt_rd_data_bits_15_11(load_io_wgt_rd_data_bits_15_11),
    .io_wgt_rd_data_bits_15_12(load_io_wgt_rd_data_bits_15_12),
    .io_wgt_rd_data_bits_15_13(load_io_wgt_rd_data_bits_15_13),
    .io_wgt_rd_data_bits_15_14(load_io_wgt_rd_data_bits_15_14),
    .io_wgt_rd_data_bits_15_15(load_io_wgt_rd_data_bits_15_15)
  );
  Compute compute ( // @[Core.scala 68:23:@24317.4]
    .clock(compute_clock),
    .reset(compute_reset),
    .io_i_post_0(compute_io_i_post_0),
    .io_i_post_1(compute_io_i_post_1),
    .io_o_post_0(compute_io_o_post_0),
    .io_o_post_1(compute_io_o_post_1),
    .io_inst_ready(compute_io_inst_ready),
    .io_inst_valid(compute_io_inst_valid),
    .io_inst_bits(compute_io_inst_bits),
    .io_uop_baddr(compute_io_uop_baddr),
    .io_acc_baddr(compute_io_acc_baddr),
    .io_vme_rd_0_cmd_ready(compute_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(compute_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(compute_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(compute_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(compute_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(compute_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits(compute_io_vme_rd_0_data_bits),
    .io_vme_rd_1_cmd_ready(compute_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(compute_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(compute_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(compute_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_data_ready(compute_io_vme_rd_1_data_ready),
    .io_vme_rd_1_data_valid(compute_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits(compute_io_vme_rd_1_data_bits),
    .io_inp_rd_idx_valid(compute_io_inp_rd_idx_valid),
    .io_inp_rd_idx_bits(compute_io_inp_rd_idx_bits),
    .io_inp_rd_data_valid(compute_io_inp_rd_data_valid),
    .io_inp_rd_data_bits_0_0(compute_io_inp_rd_data_bits_0_0),
    .io_inp_rd_data_bits_0_1(compute_io_inp_rd_data_bits_0_1),
    .io_inp_rd_data_bits_0_2(compute_io_inp_rd_data_bits_0_2),
    .io_inp_rd_data_bits_0_3(compute_io_inp_rd_data_bits_0_3),
    .io_inp_rd_data_bits_0_4(compute_io_inp_rd_data_bits_0_4),
    .io_inp_rd_data_bits_0_5(compute_io_inp_rd_data_bits_0_5),
    .io_inp_rd_data_bits_0_6(compute_io_inp_rd_data_bits_0_6),
    .io_inp_rd_data_bits_0_7(compute_io_inp_rd_data_bits_0_7),
    .io_inp_rd_data_bits_0_8(compute_io_inp_rd_data_bits_0_8),
    .io_inp_rd_data_bits_0_9(compute_io_inp_rd_data_bits_0_9),
    .io_inp_rd_data_bits_0_10(compute_io_inp_rd_data_bits_0_10),
    .io_inp_rd_data_bits_0_11(compute_io_inp_rd_data_bits_0_11),
    .io_inp_rd_data_bits_0_12(compute_io_inp_rd_data_bits_0_12),
    .io_inp_rd_data_bits_0_13(compute_io_inp_rd_data_bits_0_13),
    .io_inp_rd_data_bits_0_14(compute_io_inp_rd_data_bits_0_14),
    .io_inp_rd_data_bits_0_15(compute_io_inp_rd_data_bits_0_15),
    .io_wgt_rd_idx_valid(compute_io_wgt_rd_idx_valid),
    .io_wgt_rd_idx_bits(compute_io_wgt_rd_idx_bits),
    .io_wgt_rd_data_valid(compute_io_wgt_rd_data_valid),
    .io_wgt_rd_data_bits_0_0(compute_io_wgt_rd_data_bits_0_0),
    .io_wgt_rd_data_bits_0_1(compute_io_wgt_rd_data_bits_0_1),
    .io_wgt_rd_data_bits_0_2(compute_io_wgt_rd_data_bits_0_2),
    .io_wgt_rd_data_bits_0_3(compute_io_wgt_rd_data_bits_0_3),
    .io_wgt_rd_data_bits_0_4(compute_io_wgt_rd_data_bits_0_4),
    .io_wgt_rd_data_bits_0_5(compute_io_wgt_rd_data_bits_0_5),
    .io_wgt_rd_data_bits_0_6(compute_io_wgt_rd_data_bits_0_6),
    .io_wgt_rd_data_bits_0_7(compute_io_wgt_rd_data_bits_0_7),
    .io_wgt_rd_data_bits_0_8(compute_io_wgt_rd_data_bits_0_8),
    .io_wgt_rd_data_bits_0_9(compute_io_wgt_rd_data_bits_0_9),
    .io_wgt_rd_data_bits_0_10(compute_io_wgt_rd_data_bits_0_10),
    .io_wgt_rd_data_bits_0_11(compute_io_wgt_rd_data_bits_0_11),
    .io_wgt_rd_data_bits_0_12(compute_io_wgt_rd_data_bits_0_12),
    .io_wgt_rd_data_bits_0_13(compute_io_wgt_rd_data_bits_0_13),
    .io_wgt_rd_data_bits_0_14(compute_io_wgt_rd_data_bits_0_14),
    .io_wgt_rd_data_bits_0_15(compute_io_wgt_rd_data_bits_0_15),
    .io_wgt_rd_data_bits_1_0(compute_io_wgt_rd_data_bits_1_0),
    .io_wgt_rd_data_bits_1_1(compute_io_wgt_rd_data_bits_1_1),
    .io_wgt_rd_data_bits_1_2(compute_io_wgt_rd_data_bits_1_2),
    .io_wgt_rd_data_bits_1_3(compute_io_wgt_rd_data_bits_1_3),
    .io_wgt_rd_data_bits_1_4(compute_io_wgt_rd_data_bits_1_4),
    .io_wgt_rd_data_bits_1_5(compute_io_wgt_rd_data_bits_1_5),
    .io_wgt_rd_data_bits_1_6(compute_io_wgt_rd_data_bits_1_6),
    .io_wgt_rd_data_bits_1_7(compute_io_wgt_rd_data_bits_1_7),
    .io_wgt_rd_data_bits_1_8(compute_io_wgt_rd_data_bits_1_8),
    .io_wgt_rd_data_bits_1_9(compute_io_wgt_rd_data_bits_1_9),
    .io_wgt_rd_data_bits_1_10(compute_io_wgt_rd_data_bits_1_10),
    .io_wgt_rd_data_bits_1_11(compute_io_wgt_rd_data_bits_1_11),
    .io_wgt_rd_data_bits_1_12(compute_io_wgt_rd_data_bits_1_12),
    .io_wgt_rd_data_bits_1_13(compute_io_wgt_rd_data_bits_1_13),
    .io_wgt_rd_data_bits_1_14(compute_io_wgt_rd_data_bits_1_14),
    .io_wgt_rd_data_bits_1_15(compute_io_wgt_rd_data_bits_1_15),
    .io_wgt_rd_data_bits_2_0(compute_io_wgt_rd_data_bits_2_0),
    .io_wgt_rd_data_bits_2_1(compute_io_wgt_rd_data_bits_2_1),
    .io_wgt_rd_data_bits_2_2(compute_io_wgt_rd_data_bits_2_2),
    .io_wgt_rd_data_bits_2_3(compute_io_wgt_rd_data_bits_2_3),
    .io_wgt_rd_data_bits_2_4(compute_io_wgt_rd_data_bits_2_4),
    .io_wgt_rd_data_bits_2_5(compute_io_wgt_rd_data_bits_2_5),
    .io_wgt_rd_data_bits_2_6(compute_io_wgt_rd_data_bits_2_6),
    .io_wgt_rd_data_bits_2_7(compute_io_wgt_rd_data_bits_2_7),
    .io_wgt_rd_data_bits_2_8(compute_io_wgt_rd_data_bits_2_8),
    .io_wgt_rd_data_bits_2_9(compute_io_wgt_rd_data_bits_2_9),
    .io_wgt_rd_data_bits_2_10(compute_io_wgt_rd_data_bits_2_10),
    .io_wgt_rd_data_bits_2_11(compute_io_wgt_rd_data_bits_2_11),
    .io_wgt_rd_data_bits_2_12(compute_io_wgt_rd_data_bits_2_12),
    .io_wgt_rd_data_bits_2_13(compute_io_wgt_rd_data_bits_2_13),
    .io_wgt_rd_data_bits_2_14(compute_io_wgt_rd_data_bits_2_14),
    .io_wgt_rd_data_bits_2_15(compute_io_wgt_rd_data_bits_2_15),
    .io_wgt_rd_data_bits_3_0(compute_io_wgt_rd_data_bits_3_0),
    .io_wgt_rd_data_bits_3_1(compute_io_wgt_rd_data_bits_3_1),
    .io_wgt_rd_data_bits_3_2(compute_io_wgt_rd_data_bits_3_2),
    .io_wgt_rd_data_bits_3_3(compute_io_wgt_rd_data_bits_3_3),
    .io_wgt_rd_data_bits_3_4(compute_io_wgt_rd_data_bits_3_4),
    .io_wgt_rd_data_bits_3_5(compute_io_wgt_rd_data_bits_3_5),
    .io_wgt_rd_data_bits_3_6(compute_io_wgt_rd_data_bits_3_6),
    .io_wgt_rd_data_bits_3_7(compute_io_wgt_rd_data_bits_3_7),
    .io_wgt_rd_data_bits_3_8(compute_io_wgt_rd_data_bits_3_8),
    .io_wgt_rd_data_bits_3_9(compute_io_wgt_rd_data_bits_3_9),
    .io_wgt_rd_data_bits_3_10(compute_io_wgt_rd_data_bits_3_10),
    .io_wgt_rd_data_bits_3_11(compute_io_wgt_rd_data_bits_3_11),
    .io_wgt_rd_data_bits_3_12(compute_io_wgt_rd_data_bits_3_12),
    .io_wgt_rd_data_bits_3_13(compute_io_wgt_rd_data_bits_3_13),
    .io_wgt_rd_data_bits_3_14(compute_io_wgt_rd_data_bits_3_14),
    .io_wgt_rd_data_bits_3_15(compute_io_wgt_rd_data_bits_3_15),
    .io_wgt_rd_data_bits_4_0(compute_io_wgt_rd_data_bits_4_0),
    .io_wgt_rd_data_bits_4_1(compute_io_wgt_rd_data_bits_4_1),
    .io_wgt_rd_data_bits_4_2(compute_io_wgt_rd_data_bits_4_2),
    .io_wgt_rd_data_bits_4_3(compute_io_wgt_rd_data_bits_4_3),
    .io_wgt_rd_data_bits_4_4(compute_io_wgt_rd_data_bits_4_4),
    .io_wgt_rd_data_bits_4_5(compute_io_wgt_rd_data_bits_4_5),
    .io_wgt_rd_data_bits_4_6(compute_io_wgt_rd_data_bits_4_6),
    .io_wgt_rd_data_bits_4_7(compute_io_wgt_rd_data_bits_4_7),
    .io_wgt_rd_data_bits_4_8(compute_io_wgt_rd_data_bits_4_8),
    .io_wgt_rd_data_bits_4_9(compute_io_wgt_rd_data_bits_4_9),
    .io_wgt_rd_data_bits_4_10(compute_io_wgt_rd_data_bits_4_10),
    .io_wgt_rd_data_bits_4_11(compute_io_wgt_rd_data_bits_4_11),
    .io_wgt_rd_data_bits_4_12(compute_io_wgt_rd_data_bits_4_12),
    .io_wgt_rd_data_bits_4_13(compute_io_wgt_rd_data_bits_4_13),
    .io_wgt_rd_data_bits_4_14(compute_io_wgt_rd_data_bits_4_14),
    .io_wgt_rd_data_bits_4_15(compute_io_wgt_rd_data_bits_4_15),
    .io_wgt_rd_data_bits_5_0(compute_io_wgt_rd_data_bits_5_0),
    .io_wgt_rd_data_bits_5_1(compute_io_wgt_rd_data_bits_5_1),
    .io_wgt_rd_data_bits_5_2(compute_io_wgt_rd_data_bits_5_2),
    .io_wgt_rd_data_bits_5_3(compute_io_wgt_rd_data_bits_5_3),
    .io_wgt_rd_data_bits_5_4(compute_io_wgt_rd_data_bits_5_4),
    .io_wgt_rd_data_bits_5_5(compute_io_wgt_rd_data_bits_5_5),
    .io_wgt_rd_data_bits_5_6(compute_io_wgt_rd_data_bits_5_6),
    .io_wgt_rd_data_bits_5_7(compute_io_wgt_rd_data_bits_5_7),
    .io_wgt_rd_data_bits_5_8(compute_io_wgt_rd_data_bits_5_8),
    .io_wgt_rd_data_bits_5_9(compute_io_wgt_rd_data_bits_5_9),
    .io_wgt_rd_data_bits_5_10(compute_io_wgt_rd_data_bits_5_10),
    .io_wgt_rd_data_bits_5_11(compute_io_wgt_rd_data_bits_5_11),
    .io_wgt_rd_data_bits_5_12(compute_io_wgt_rd_data_bits_5_12),
    .io_wgt_rd_data_bits_5_13(compute_io_wgt_rd_data_bits_5_13),
    .io_wgt_rd_data_bits_5_14(compute_io_wgt_rd_data_bits_5_14),
    .io_wgt_rd_data_bits_5_15(compute_io_wgt_rd_data_bits_5_15),
    .io_wgt_rd_data_bits_6_0(compute_io_wgt_rd_data_bits_6_0),
    .io_wgt_rd_data_bits_6_1(compute_io_wgt_rd_data_bits_6_1),
    .io_wgt_rd_data_bits_6_2(compute_io_wgt_rd_data_bits_6_2),
    .io_wgt_rd_data_bits_6_3(compute_io_wgt_rd_data_bits_6_3),
    .io_wgt_rd_data_bits_6_4(compute_io_wgt_rd_data_bits_6_4),
    .io_wgt_rd_data_bits_6_5(compute_io_wgt_rd_data_bits_6_5),
    .io_wgt_rd_data_bits_6_6(compute_io_wgt_rd_data_bits_6_6),
    .io_wgt_rd_data_bits_6_7(compute_io_wgt_rd_data_bits_6_7),
    .io_wgt_rd_data_bits_6_8(compute_io_wgt_rd_data_bits_6_8),
    .io_wgt_rd_data_bits_6_9(compute_io_wgt_rd_data_bits_6_9),
    .io_wgt_rd_data_bits_6_10(compute_io_wgt_rd_data_bits_6_10),
    .io_wgt_rd_data_bits_6_11(compute_io_wgt_rd_data_bits_6_11),
    .io_wgt_rd_data_bits_6_12(compute_io_wgt_rd_data_bits_6_12),
    .io_wgt_rd_data_bits_6_13(compute_io_wgt_rd_data_bits_6_13),
    .io_wgt_rd_data_bits_6_14(compute_io_wgt_rd_data_bits_6_14),
    .io_wgt_rd_data_bits_6_15(compute_io_wgt_rd_data_bits_6_15),
    .io_wgt_rd_data_bits_7_0(compute_io_wgt_rd_data_bits_7_0),
    .io_wgt_rd_data_bits_7_1(compute_io_wgt_rd_data_bits_7_1),
    .io_wgt_rd_data_bits_7_2(compute_io_wgt_rd_data_bits_7_2),
    .io_wgt_rd_data_bits_7_3(compute_io_wgt_rd_data_bits_7_3),
    .io_wgt_rd_data_bits_7_4(compute_io_wgt_rd_data_bits_7_4),
    .io_wgt_rd_data_bits_7_5(compute_io_wgt_rd_data_bits_7_5),
    .io_wgt_rd_data_bits_7_6(compute_io_wgt_rd_data_bits_7_6),
    .io_wgt_rd_data_bits_7_7(compute_io_wgt_rd_data_bits_7_7),
    .io_wgt_rd_data_bits_7_8(compute_io_wgt_rd_data_bits_7_8),
    .io_wgt_rd_data_bits_7_9(compute_io_wgt_rd_data_bits_7_9),
    .io_wgt_rd_data_bits_7_10(compute_io_wgt_rd_data_bits_7_10),
    .io_wgt_rd_data_bits_7_11(compute_io_wgt_rd_data_bits_7_11),
    .io_wgt_rd_data_bits_7_12(compute_io_wgt_rd_data_bits_7_12),
    .io_wgt_rd_data_bits_7_13(compute_io_wgt_rd_data_bits_7_13),
    .io_wgt_rd_data_bits_7_14(compute_io_wgt_rd_data_bits_7_14),
    .io_wgt_rd_data_bits_7_15(compute_io_wgt_rd_data_bits_7_15),
    .io_wgt_rd_data_bits_8_0(compute_io_wgt_rd_data_bits_8_0),
    .io_wgt_rd_data_bits_8_1(compute_io_wgt_rd_data_bits_8_1),
    .io_wgt_rd_data_bits_8_2(compute_io_wgt_rd_data_bits_8_2),
    .io_wgt_rd_data_bits_8_3(compute_io_wgt_rd_data_bits_8_3),
    .io_wgt_rd_data_bits_8_4(compute_io_wgt_rd_data_bits_8_4),
    .io_wgt_rd_data_bits_8_5(compute_io_wgt_rd_data_bits_8_5),
    .io_wgt_rd_data_bits_8_6(compute_io_wgt_rd_data_bits_8_6),
    .io_wgt_rd_data_bits_8_7(compute_io_wgt_rd_data_bits_8_7),
    .io_wgt_rd_data_bits_8_8(compute_io_wgt_rd_data_bits_8_8),
    .io_wgt_rd_data_bits_8_9(compute_io_wgt_rd_data_bits_8_9),
    .io_wgt_rd_data_bits_8_10(compute_io_wgt_rd_data_bits_8_10),
    .io_wgt_rd_data_bits_8_11(compute_io_wgt_rd_data_bits_8_11),
    .io_wgt_rd_data_bits_8_12(compute_io_wgt_rd_data_bits_8_12),
    .io_wgt_rd_data_bits_8_13(compute_io_wgt_rd_data_bits_8_13),
    .io_wgt_rd_data_bits_8_14(compute_io_wgt_rd_data_bits_8_14),
    .io_wgt_rd_data_bits_8_15(compute_io_wgt_rd_data_bits_8_15),
    .io_wgt_rd_data_bits_9_0(compute_io_wgt_rd_data_bits_9_0),
    .io_wgt_rd_data_bits_9_1(compute_io_wgt_rd_data_bits_9_1),
    .io_wgt_rd_data_bits_9_2(compute_io_wgt_rd_data_bits_9_2),
    .io_wgt_rd_data_bits_9_3(compute_io_wgt_rd_data_bits_9_3),
    .io_wgt_rd_data_bits_9_4(compute_io_wgt_rd_data_bits_9_4),
    .io_wgt_rd_data_bits_9_5(compute_io_wgt_rd_data_bits_9_5),
    .io_wgt_rd_data_bits_9_6(compute_io_wgt_rd_data_bits_9_6),
    .io_wgt_rd_data_bits_9_7(compute_io_wgt_rd_data_bits_9_7),
    .io_wgt_rd_data_bits_9_8(compute_io_wgt_rd_data_bits_9_8),
    .io_wgt_rd_data_bits_9_9(compute_io_wgt_rd_data_bits_9_9),
    .io_wgt_rd_data_bits_9_10(compute_io_wgt_rd_data_bits_9_10),
    .io_wgt_rd_data_bits_9_11(compute_io_wgt_rd_data_bits_9_11),
    .io_wgt_rd_data_bits_9_12(compute_io_wgt_rd_data_bits_9_12),
    .io_wgt_rd_data_bits_9_13(compute_io_wgt_rd_data_bits_9_13),
    .io_wgt_rd_data_bits_9_14(compute_io_wgt_rd_data_bits_9_14),
    .io_wgt_rd_data_bits_9_15(compute_io_wgt_rd_data_bits_9_15),
    .io_wgt_rd_data_bits_10_0(compute_io_wgt_rd_data_bits_10_0),
    .io_wgt_rd_data_bits_10_1(compute_io_wgt_rd_data_bits_10_1),
    .io_wgt_rd_data_bits_10_2(compute_io_wgt_rd_data_bits_10_2),
    .io_wgt_rd_data_bits_10_3(compute_io_wgt_rd_data_bits_10_3),
    .io_wgt_rd_data_bits_10_4(compute_io_wgt_rd_data_bits_10_4),
    .io_wgt_rd_data_bits_10_5(compute_io_wgt_rd_data_bits_10_5),
    .io_wgt_rd_data_bits_10_6(compute_io_wgt_rd_data_bits_10_6),
    .io_wgt_rd_data_bits_10_7(compute_io_wgt_rd_data_bits_10_7),
    .io_wgt_rd_data_bits_10_8(compute_io_wgt_rd_data_bits_10_8),
    .io_wgt_rd_data_bits_10_9(compute_io_wgt_rd_data_bits_10_9),
    .io_wgt_rd_data_bits_10_10(compute_io_wgt_rd_data_bits_10_10),
    .io_wgt_rd_data_bits_10_11(compute_io_wgt_rd_data_bits_10_11),
    .io_wgt_rd_data_bits_10_12(compute_io_wgt_rd_data_bits_10_12),
    .io_wgt_rd_data_bits_10_13(compute_io_wgt_rd_data_bits_10_13),
    .io_wgt_rd_data_bits_10_14(compute_io_wgt_rd_data_bits_10_14),
    .io_wgt_rd_data_bits_10_15(compute_io_wgt_rd_data_bits_10_15),
    .io_wgt_rd_data_bits_11_0(compute_io_wgt_rd_data_bits_11_0),
    .io_wgt_rd_data_bits_11_1(compute_io_wgt_rd_data_bits_11_1),
    .io_wgt_rd_data_bits_11_2(compute_io_wgt_rd_data_bits_11_2),
    .io_wgt_rd_data_bits_11_3(compute_io_wgt_rd_data_bits_11_3),
    .io_wgt_rd_data_bits_11_4(compute_io_wgt_rd_data_bits_11_4),
    .io_wgt_rd_data_bits_11_5(compute_io_wgt_rd_data_bits_11_5),
    .io_wgt_rd_data_bits_11_6(compute_io_wgt_rd_data_bits_11_6),
    .io_wgt_rd_data_bits_11_7(compute_io_wgt_rd_data_bits_11_7),
    .io_wgt_rd_data_bits_11_8(compute_io_wgt_rd_data_bits_11_8),
    .io_wgt_rd_data_bits_11_9(compute_io_wgt_rd_data_bits_11_9),
    .io_wgt_rd_data_bits_11_10(compute_io_wgt_rd_data_bits_11_10),
    .io_wgt_rd_data_bits_11_11(compute_io_wgt_rd_data_bits_11_11),
    .io_wgt_rd_data_bits_11_12(compute_io_wgt_rd_data_bits_11_12),
    .io_wgt_rd_data_bits_11_13(compute_io_wgt_rd_data_bits_11_13),
    .io_wgt_rd_data_bits_11_14(compute_io_wgt_rd_data_bits_11_14),
    .io_wgt_rd_data_bits_11_15(compute_io_wgt_rd_data_bits_11_15),
    .io_wgt_rd_data_bits_12_0(compute_io_wgt_rd_data_bits_12_0),
    .io_wgt_rd_data_bits_12_1(compute_io_wgt_rd_data_bits_12_1),
    .io_wgt_rd_data_bits_12_2(compute_io_wgt_rd_data_bits_12_2),
    .io_wgt_rd_data_bits_12_3(compute_io_wgt_rd_data_bits_12_3),
    .io_wgt_rd_data_bits_12_4(compute_io_wgt_rd_data_bits_12_4),
    .io_wgt_rd_data_bits_12_5(compute_io_wgt_rd_data_bits_12_5),
    .io_wgt_rd_data_bits_12_6(compute_io_wgt_rd_data_bits_12_6),
    .io_wgt_rd_data_bits_12_7(compute_io_wgt_rd_data_bits_12_7),
    .io_wgt_rd_data_bits_12_8(compute_io_wgt_rd_data_bits_12_8),
    .io_wgt_rd_data_bits_12_9(compute_io_wgt_rd_data_bits_12_9),
    .io_wgt_rd_data_bits_12_10(compute_io_wgt_rd_data_bits_12_10),
    .io_wgt_rd_data_bits_12_11(compute_io_wgt_rd_data_bits_12_11),
    .io_wgt_rd_data_bits_12_12(compute_io_wgt_rd_data_bits_12_12),
    .io_wgt_rd_data_bits_12_13(compute_io_wgt_rd_data_bits_12_13),
    .io_wgt_rd_data_bits_12_14(compute_io_wgt_rd_data_bits_12_14),
    .io_wgt_rd_data_bits_12_15(compute_io_wgt_rd_data_bits_12_15),
    .io_wgt_rd_data_bits_13_0(compute_io_wgt_rd_data_bits_13_0),
    .io_wgt_rd_data_bits_13_1(compute_io_wgt_rd_data_bits_13_1),
    .io_wgt_rd_data_bits_13_2(compute_io_wgt_rd_data_bits_13_2),
    .io_wgt_rd_data_bits_13_3(compute_io_wgt_rd_data_bits_13_3),
    .io_wgt_rd_data_bits_13_4(compute_io_wgt_rd_data_bits_13_4),
    .io_wgt_rd_data_bits_13_5(compute_io_wgt_rd_data_bits_13_5),
    .io_wgt_rd_data_bits_13_6(compute_io_wgt_rd_data_bits_13_6),
    .io_wgt_rd_data_bits_13_7(compute_io_wgt_rd_data_bits_13_7),
    .io_wgt_rd_data_bits_13_8(compute_io_wgt_rd_data_bits_13_8),
    .io_wgt_rd_data_bits_13_9(compute_io_wgt_rd_data_bits_13_9),
    .io_wgt_rd_data_bits_13_10(compute_io_wgt_rd_data_bits_13_10),
    .io_wgt_rd_data_bits_13_11(compute_io_wgt_rd_data_bits_13_11),
    .io_wgt_rd_data_bits_13_12(compute_io_wgt_rd_data_bits_13_12),
    .io_wgt_rd_data_bits_13_13(compute_io_wgt_rd_data_bits_13_13),
    .io_wgt_rd_data_bits_13_14(compute_io_wgt_rd_data_bits_13_14),
    .io_wgt_rd_data_bits_13_15(compute_io_wgt_rd_data_bits_13_15),
    .io_wgt_rd_data_bits_14_0(compute_io_wgt_rd_data_bits_14_0),
    .io_wgt_rd_data_bits_14_1(compute_io_wgt_rd_data_bits_14_1),
    .io_wgt_rd_data_bits_14_2(compute_io_wgt_rd_data_bits_14_2),
    .io_wgt_rd_data_bits_14_3(compute_io_wgt_rd_data_bits_14_3),
    .io_wgt_rd_data_bits_14_4(compute_io_wgt_rd_data_bits_14_4),
    .io_wgt_rd_data_bits_14_5(compute_io_wgt_rd_data_bits_14_5),
    .io_wgt_rd_data_bits_14_6(compute_io_wgt_rd_data_bits_14_6),
    .io_wgt_rd_data_bits_14_7(compute_io_wgt_rd_data_bits_14_7),
    .io_wgt_rd_data_bits_14_8(compute_io_wgt_rd_data_bits_14_8),
    .io_wgt_rd_data_bits_14_9(compute_io_wgt_rd_data_bits_14_9),
    .io_wgt_rd_data_bits_14_10(compute_io_wgt_rd_data_bits_14_10),
    .io_wgt_rd_data_bits_14_11(compute_io_wgt_rd_data_bits_14_11),
    .io_wgt_rd_data_bits_14_12(compute_io_wgt_rd_data_bits_14_12),
    .io_wgt_rd_data_bits_14_13(compute_io_wgt_rd_data_bits_14_13),
    .io_wgt_rd_data_bits_14_14(compute_io_wgt_rd_data_bits_14_14),
    .io_wgt_rd_data_bits_14_15(compute_io_wgt_rd_data_bits_14_15),
    .io_wgt_rd_data_bits_15_0(compute_io_wgt_rd_data_bits_15_0),
    .io_wgt_rd_data_bits_15_1(compute_io_wgt_rd_data_bits_15_1),
    .io_wgt_rd_data_bits_15_2(compute_io_wgt_rd_data_bits_15_2),
    .io_wgt_rd_data_bits_15_3(compute_io_wgt_rd_data_bits_15_3),
    .io_wgt_rd_data_bits_15_4(compute_io_wgt_rd_data_bits_15_4),
    .io_wgt_rd_data_bits_15_5(compute_io_wgt_rd_data_bits_15_5),
    .io_wgt_rd_data_bits_15_6(compute_io_wgt_rd_data_bits_15_6),
    .io_wgt_rd_data_bits_15_7(compute_io_wgt_rd_data_bits_15_7),
    .io_wgt_rd_data_bits_15_8(compute_io_wgt_rd_data_bits_15_8),
    .io_wgt_rd_data_bits_15_9(compute_io_wgt_rd_data_bits_15_9),
    .io_wgt_rd_data_bits_15_10(compute_io_wgt_rd_data_bits_15_10),
    .io_wgt_rd_data_bits_15_11(compute_io_wgt_rd_data_bits_15_11),
    .io_wgt_rd_data_bits_15_12(compute_io_wgt_rd_data_bits_15_12),
    .io_wgt_rd_data_bits_15_13(compute_io_wgt_rd_data_bits_15_13),
    .io_wgt_rd_data_bits_15_14(compute_io_wgt_rd_data_bits_15_14),
    .io_wgt_rd_data_bits_15_15(compute_io_wgt_rd_data_bits_15_15),
    .io_out_wr_valid(compute_io_out_wr_valid),
    .io_out_wr_bits_idx(compute_io_out_wr_bits_idx),
    .io_out_wr_bits_data_0_0(compute_io_out_wr_bits_data_0_0),
    .io_out_wr_bits_data_0_1(compute_io_out_wr_bits_data_0_1),
    .io_out_wr_bits_data_0_2(compute_io_out_wr_bits_data_0_2),
    .io_out_wr_bits_data_0_3(compute_io_out_wr_bits_data_0_3),
    .io_out_wr_bits_data_0_4(compute_io_out_wr_bits_data_0_4),
    .io_out_wr_bits_data_0_5(compute_io_out_wr_bits_data_0_5),
    .io_out_wr_bits_data_0_6(compute_io_out_wr_bits_data_0_6),
    .io_out_wr_bits_data_0_7(compute_io_out_wr_bits_data_0_7),
    .io_out_wr_bits_data_0_8(compute_io_out_wr_bits_data_0_8),
    .io_out_wr_bits_data_0_9(compute_io_out_wr_bits_data_0_9),
    .io_out_wr_bits_data_0_10(compute_io_out_wr_bits_data_0_10),
    .io_out_wr_bits_data_0_11(compute_io_out_wr_bits_data_0_11),
    .io_out_wr_bits_data_0_12(compute_io_out_wr_bits_data_0_12),
    .io_out_wr_bits_data_0_13(compute_io_out_wr_bits_data_0_13),
    .io_out_wr_bits_data_0_14(compute_io_out_wr_bits_data_0_14),
    .io_out_wr_bits_data_0_15(compute_io_out_wr_bits_data_0_15),
    .io_finish(compute_io_finish),
    .io_acc_wr_event(compute_io_acc_wr_event)
  );
  Store store ( // @[Core.scala 69:21:@24320.4]
    .clock(store_clock),
    .reset(store_reset),
    .io_i_post(store_io_i_post),
    .io_o_post(store_io_o_post),
    .io_inst_ready(store_io_inst_ready),
    .io_inst_valid(store_io_inst_valid),
    .io_inst_bits(store_io_inst_bits),
    .io_out_baddr(store_io_out_baddr),
    .io_vme_wr_cmd_ready(store_io_vme_wr_cmd_ready),
    .io_vme_wr_cmd_valid(store_io_vme_wr_cmd_valid),
    .io_vme_wr_cmd_bits_addr(store_io_vme_wr_cmd_bits_addr),
    .io_vme_wr_cmd_bits_len(store_io_vme_wr_cmd_bits_len),
    .io_vme_wr_data_ready(store_io_vme_wr_data_ready),
    .io_vme_wr_data_valid(store_io_vme_wr_data_valid),
    .io_vme_wr_data_bits(store_io_vme_wr_data_bits),
    .io_vme_wr_ack(store_io_vme_wr_ack),
    .io_out_wr_valid(store_io_out_wr_valid),
    .io_out_wr_bits_idx(store_io_out_wr_bits_idx),
    .io_out_wr_bits_data_0_0(store_io_out_wr_bits_data_0_0),
    .io_out_wr_bits_data_0_1(store_io_out_wr_bits_data_0_1),
    .io_out_wr_bits_data_0_2(store_io_out_wr_bits_data_0_2),
    .io_out_wr_bits_data_0_3(store_io_out_wr_bits_data_0_3),
    .io_out_wr_bits_data_0_4(store_io_out_wr_bits_data_0_4),
    .io_out_wr_bits_data_0_5(store_io_out_wr_bits_data_0_5),
    .io_out_wr_bits_data_0_6(store_io_out_wr_bits_data_0_6),
    .io_out_wr_bits_data_0_7(store_io_out_wr_bits_data_0_7),
    .io_out_wr_bits_data_0_8(store_io_out_wr_bits_data_0_8),
    .io_out_wr_bits_data_0_9(store_io_out_wr_bits_data_0_9),
    .io_out_wr_bits_data_0_10(store_io_out_wr_bits_data_0_10),
    .io_out_wr_bits_data_0_11(store_io_out_wr_bits_data_0_11),
    .io_out_wr_bits_data_0_12(store_io_out_wr_bits_data_0_12),
    .io_out_wr_bits_data_0_13(store_io_out_wr_bits_data_0_13),
    .io_out_wr_bits_data_0_14(store_io_out_wr_bits_data_0_14),
    .io_out_wr_bits_data_0_15(store_io_out_wr_bits_data_0_15)
  );
  EventCounters ecounters ( // @[Core.scala 70:25:@24323.4]
    .clock(ecounters_clock),
    .reset(ecounters_reset),
    .io_launch(ecounters_io_launch),
    .io_finish(ecounters_io_finish),
    .io_ecnt_0_valid(ecounters_io_ecnt_0_valid),
    .io_ecnt_0_bits(ecounters_io_ecnt_0_bits),
    .io_ucnt_0_valid(ecounters_io_ucnt_0_valid),
    .io_ucnt_0_bits(ecounters_io_ucnt_0_bits),
    .io_acc_wr_event(ecounters_io_acc_wr_event)
  );
  assign io_vcr_finish = finish; // @[Core.scala 119:17:@24990.4]
  assign io_vcr_ecnt_0_valid = ecounters_io_ecnt_0_valid; // @[Core.scala 113:15:@24984.4]
  assign io_vcr_ecnt_0_bits = ecounters_io_ecnt_0_bits; // @[Core.scala 113:15:@24983.4]
  assign io_vcr_ucnt_0_valid = ecounters_io_ucnt_0_valid; // @[Core.scala 114:15:@24986.4]
  assign io_vcr_ucnt_0_bits = ecounters_io_ucnt_0_bits; // @[Core.scala 114:15:@24985.4]
  assign io_vme_rd_0_cmd_valid = fetch_io_vme_rd_cmd_valid; // @[Core.scala 73:16:@24331.4]
  assign io_vme_rd_0_cmd_bits_addr = fetch_io_vme_rd_cmd_bits_addr; // @[Core.scala 73:16:@24330.4]
  assign io_vme_rd_0_cmd_bits_len = fetch_io_vme_rd_cmd_bits_len; // @[Core.scala 73:16:@24329.4]
  assign io_vme_rd_0_data_ready = fetch_io_vme_rd_data_ready; // @[Core.scala 73:16:@24328.4]
  assign io_vme_rd_1_cmd_valid = compute_io_vme_rd_0_cmd_valid; // @[Core.scala 74:16:@24338.4]
  assign io_vme_rd_1_cmd_bits_addr = compute_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 74:16:@24337.4]
  assign io_vme_rd_1_cmd_bits_len = compute_io_vme_rd_0_cmd_bits_len; // @[Core.scala 74:16:@24336.4]
  assign io_vme_rd_1_data_ready = compute_io_vme_rd_0_data_ready; // @[Core.scala 74:16:@24335.4]
  assign io_vme_rd_2_cmd_valid = load_io_vme_rd_0_cmd_valid; // @[Core.scala 75:16:@24345.4]
  assign io_vme_rd_2_cmd_bits_addr = load_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 75:16:@24344.4]
  assign io_vme_rd_2_cmd_bits_len = load_io_vme_rd_0_cmd_bits_len; // @[Core.scala 75:16:@24343.4]
  assign io_vme_rd_2_data_ready = load_io_vme_rd_0_data_ready; // @[Core.scala 75:16:@24342.4]
  assign io_vme_rd_3_cmd_valid = load_io_vme_rd_1_cmd_valid; // @[Core.scala 76:16:@24352.4]
  assign io_vme_rd_3_cmd_bits_addr = load_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 76:16:@24351.4]
  assign io_vme_rd_3_cmd_bits_len = load_io_vme_rd_1_cmd_bits_len; // @[Core.scala 76:16:@24350.4]
  assign io_vme_rd_3_data_ready = load_io_vme_rd_1_data_ready; // @[Core.scala 76:16:@24349.4]
  assign io_vme_rd_4_cmd_valid = compute_io_vme_rd_1_cmd_valid; // @[Core.scala 77:16:@24359.4]
  assign io_vme_rd_4_cmd_bits_addr = compute_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 77:16:@24358.4]
  assign io_vme_rd_4_cmd_bits_len = compute_io_vme_rd_1_cmd_bits_len; // @[Core.scala 77:16:@24357.4]
  assign io_vme_rd_4_data_ready = compute_io_vme_rd_1_data_ready; // @[Core.scala 77:16:@24356.4]
  assign io_vme_wr_0_cmd_valid = store_io_vme_wr_cmd_valid; // @[Core.scala 78:16:@24367.4]
  assign io_vme_wr_0_cmd_bits_addr = store_io_vme_wr_cmd_bits_addr; // @[Core.scala 78:16:@24366.4]
  assign io_vme_wr_0_cmd_bits_len = store_io_vme_wr_cmd_bits_len; // @[Core.scala 78:16:@24365.4]
  assign io_vme_wr_0_data_valid = store_io_vme_wr_data_valid; // @[Core.scala 78:16:@24363.4]
  assign io_vme_wr_0_data_bits = store_io_vme_wr_data_bits; // @[Core.scala 78:16:@24362.4]
  assign fetch_clock = clock; // @[:@24312.4]
  assign fetch_reset = reset; // @[:@24313.4]
  assign fetch_io_launch = io_vcr_launch; // @[Core.scala 81:19:@24369.4]
  assign fetch_io_ins_baddr = io_vcr_ptrs_0; // @[Core.scala 82:22:@24370.4]
  assign fetch_io_ins_count = io_vcr_vals_0; // @[Core.scala 83:22:@24371.4]
  assign fetch_io_vme_rd_cmd_ready = io_vme_rd_0_cmd_ready; // @[Core.scala 73:16:@24332.4]
  assign fetch_io_vme_rd_data_valid = io_vme_rd_0_data_valid; // @[Core.scala 73:16:@24327.4]
  assign fetch_io_vme_rd_data_bits = io_vme_rd_0_data_bits; // @[Core.scala 73:16:@24326.4]
  assign fetch_io_inst_ld_ready = load_io_inst_ready; // @[Core.scala 87:16:@24375.4]
  assign fetch_io_inst_co_ready = compute_io_inst_ready; // @[Core.scala 96:19:@24382.4]
  assign fetch_io_inst_st_ready = store_io_inst_ready; // @[Core.scala 106:17:@24942.4]
  assign load_clock = clock; // @[:@24315.4]
  assign load_reset = reset; // @[:@24316.4]
  assign load_io_i_post = compute_io_o_post_0; // @[Core.scala 86:18:@24372.4]
  assign load_io_inst_valid = fetch_io_inst_ld_valid; // @[Core.scala 87:16:@24374.4]
  assign load_io_inst_bits = fetch_io_inst_ld_bits; // @[Core.scala 87:16:@24373.4]
  assign load_io_inp_baddr = io_vcr_ptrs_2; // @[Core.scala 88:21:@24376.4]
  assign load_io_wgt_baddr = io_vcr_ptrs_3; // @[Core.scala 89:21:@24377.4]
  assign load_io_vme_rd_0_cmd_ready = io_vme_rd_2_cmd_ready; // @[Core.scala 75:16:@24346.4]
  assign load_io_vme_rd_0_data_valid = io_vme_rd_2_data_valid; // @[Core.scala 75:16:@24341.4]
  assign load_io_vme_rd_0_data_bits = io_vme_rd_2_data_bits; // @[Core.scala 75:16:@24340.4]
  assign load_io_vme_rd_1_cmd_ready = io_vme_rd_3_cmd_ready; // @[Core.scala 76:16:@24353.4]
  assign load_io_vme_rd_1_data_valid = io_vme_rd_3_data_valid; // @[Core.scala 76:16:@24348.4]
  assign load_io_vme_rd_1_data_bits = io_vme_rd_3_data_bits; // @[Core.scala 76:16:@24347.4]
  assign load_io_inp_rd_idx_valid = compute_io_inp_rd_idx_valid; // @[Core.scala 99:18:@24421.4]
  assign load_io_inp_rd_idx_bits = compute_io_inp_rd_idx_bits; // @[Core.scala 99:18:@24420.4]
  assign load_io_wgt_rd_idx_valid = compute_io_wgt_rd_idx_valid; // @[Core.scala 100:18:@24938.4]
  assign load_io_wgt_rd_idx_bits = compute_io_wgt_rd_idx_bits; // @[Core.scala 100:18:@24937.4]
  assign compute_clock = clock; // @[:@24318.4]
  assign compute_reset = reset; // @[:@24319.4]
  assign compute_io_i_post_0 = load_io_o_post; // @[Core.scala 94:24:@24378.4]
  assign compute_io_i_post_1 = store_io_o_post; // @[Core.scala 95:24:@24379.4]
  assign compute_io_inst_valid = fetch_io_inst_co_valid; // @[Core.scala 96:19:@24381.4]
  assign compute_io_inst_bits = fetch_io_inst_co_bits; // @[Core.scala 96:19:@24380.4]
  assign compute_io_uop_baddr = io_vcr_ptrs_1; // @[Core.scala 97:24:@24383.4]
  assign compute_io_acc_baddr = io_vcr_ptrs_4; // @[Core.scala 98:24:@24384.4]
  assign compute_io_vme_rd_0_cmd_ready = io_vme_rd_1_cmd_ready; // @[Core.scala 74:16:@24339.4]
  assign compute_io_vme_rd_0_data_valid = io_vme_rd_1_data_valid; // @[Core.scala 74:16:@24334.4]
  assign compute_io_vme_rd_0_data_bits = io_vme_rd_1_data_bits; // @[Core.scala 74:16:@24333.4]
  assign compute_io_vme_rd_1_cmd_ready = io_vme_rd_4_cmd_ready; // @[Core.scala 77:16:@24360.4]
  assign compute_io_vme_rd_1_data_valid = io_vme_rd_4_data_valid; // @[Core.scala 77:16:@24355.4]
  assign compute_io_vme_rd_1_data_bits = io_vme_rd_4_data_bits; // @[Core.scala 77:16:@24354.4]
  assign compute_io_inp_rd_data_valid = load_io_inp_rd_data_valid; // @[Core.scala 99:18:@24419.4]
  assign compute_io_inp_rd_data_bits_0_0 = load_io_inp_rd_data_bits_0_0; // @[Core.scala 99:18:@24403.4]
  assign compute_io_inp_rd_data_bits_0_1 = load_io_inp_rd_data_bits_0_1; // @[Core.scala 99:18:@24404.4]
  assign compute_io_inp_rd_data_bits_0_2 = load_io_inp_rd_data_bits_0_2; // @[Core.scala 99:18:@24405.4]
  assign compute_io_inp_rd_data_bits_0_3 = load_io_inp_rd_data_bits_0_3; // @[Core.scala 99:18:@24406.4]
  assign compute_io_inp_rd_data_bits_0_4 = load_io_inp_rd_data_bits_0_4; // @[Core.scala 99:18:@24407.4]
  assign compute_io_inp_rd_data_bits_0_5 = load_io_inp_rd_data_bits_0_5; // @[Core.scala 99:18:@24408.4]
  assign compute_io_inp_rd_data_bits_0_6 = load_io_inp_rd_data_bits_0_6; // @[Core.scala 99:18:@24409.4]
  assign compute_io_inp_rd_data_bits_0_7 = load_io_inp_rd_data_bits_0_7; // @[Core.scala 99:18:@24410.4]
  assign compute_io_inp_rd_data_bits_0_8 = load_io_inp_rd_data_bits_0_8; // @[Core.scala 99:18:@24411.4]
  assign compute_io_inp_rd_data_bits_0_9 = load_io_inp_rd_data_bits_0_9; // @[Core.scala 99:18:@24412.4]
  assign compute_io_inp_rd_data_bits_0_10 = load_io_inp_rd_data_bits_0_10; // @[Core.scala 99:18:@24413.4]
  assign compute_io_inp_rd_data_bits_0_11 = load_io_inp_rd_data_bits_0_11; // @[Core.scala 99:18:@24414.4]
  assign compute_io_inp_rd_data_bits_0_12 = load_io_inp_rd_data_bits_0_12; // @[Core.scala 99:18:@24415.4]
  assign compute_io_inp_rd_data_bits_0_13 = load_io_inp_rd_data_bits_0_13; // @[Core.scala 99:18:@24416.4]
  assign compute_io_inp_rd_data_bits_0_14 = load_io_inp_rd_data_bits_0_14; // @[Core.scala 99:18:@24417.4]
  assign compute_io_inp_rd_data_bits_0_15 = load_io_inp_rd_data_bits_0_15; // @[Core.scala 99:18:@24418.4]
  assign compute_io_wgt_rd_data_valid = load_io_wgt_rd_data_valid; // @[Core.scala 100:18:@24936.4]
  assign compute_io_wgt_rd_data_bits_0_0 = load_io_wgt_rd_data_bits_0_0; // @[Core.scala 100:18:@24680.4]
  assign compute_io_wgt_rd_data_bits_0_1 = load_io_wgt_rd_data_bits_0_1; // @[Core.scala 100:18:@24681.4]
  assign compute_io_wgt_rd_data_bits_0_2 = load_io_wgt_rd_data_bits_0_2; // @[Core.scala 100:18:@24682.4]
  assign compute_io_wgt_rd_data_bits_0_3 = load_io_wgt_rd_data_bits_0_3; // @[Core.scala 100:18:@24683.4]
  assign compute_io_wgt_rd_data_bits_0_4 = load_io_wgt_rd_data_bits_0_4; // @[Core.scala 100:18:@24684.4]
  assign compute_io_wgt_rd_data_bits_0_5 = load_io_wgt_rd_data_bits_0_5; // @[Core.scala 100:18:@24685.4]
  assign compute_io_wgt_rd_data_bits_0_6 = load_io_wgt_rd_data_bits_0_6; // @[Core.scala 100:18:@24686.4]
  assign compute_io_wgt_rd_data_bits_0_7 = load_io_wgt_rd_data_bits_0_7; // @[Core.scala 100:18:@24687.4]
  assign compute_io_wgt_rd_data_bits_0_8 = load_io_wgt_rd_data_bits_0_8; // @[Core.scala 100:18:@24688.4]
  assign compute_io_wgt_rd_data_bits_0_9 = load_io_wgt_rd_data_bits_0_9; // @[Core.scala 100:18:@24689.4]
  assign compute_io_wgt_rd_data_bits_0_10 = load_io_wgt_rd_data_bits_0_10; // @[Core.scala 100:18:@24690.4]
  assign compute_io_wgt_rd_data_bits_0_11 = load_io_wgt_rd_data_bits_0_11; // @[Core.scala 100:18:@24691.4]
  assign compute_io_wgt_rd_data_bits_0_12 = load_io_wgt_rd_data_bits_0_12; // @[Core.scala 100:18:@24692.4]
  assign compute_io_wgt_rd_data_bits_0_13 = load_io_wgt_rd_data_bits_0_13; // @[Core.scala 100:18:@24693.4]
  assign compute_io_wgt_rd_data_bits_0_14 = load_io_wgt_rd_data_bits_0_14; // @[Core.scala 100:18:@24694.4]
  assign compute_io_wgt_rd_data_bits_0_15 = load_io_wgt_rd_data_bits_0_15; // @[Core.scala 100:18:@24695.4]
  assign compute_io_wgt_rd_data_bits_1_0 = load_io_wgt_rd_data_bits_1_0; // @[Core.scala 100:18:@24696.4]
  assign compute_io_wgt_rd_data_bits_1_1 = load_io_wgt_rd_data_bits_1_1; // @[Core.scala 100:18:@24697.4]
  assign compute_io_wgt_rd_data_bits_1_2 = load_io_wgt_rd_data_bits_1_2; // @[Core.scala 100:18:@24698.4]
  assign compute_io_wgt_rd_data_bits_1_3 = load_io_wgt_rd_data_bits_1_3; // @[Core.scala 100:18:@24699.4]
  assign compute_io_wgt_rd_data_bits_1_4 = load_io_wgt_rd_data_bits_1_4; // @[Core.scala 100:18:@24700.4]
  assign compute_io_wgt_rd_data_bits_1_5 = load_io_wgt_rd_data_bits_1_5; // @[Core.scala 100:18:@24701.4]
  assign compute_io_wgt_rd_data_bits_1_6 = load_io_wgt_rd_data_bits_1_6; // @[Core.scala 100:18:@24702.4]
  assign compute_io_wgt_rd_data_bits_1_7 = load_io_wgt_rd_data_bits_1_7; // @[Core.scala 100:18:@24703.4]
  assign compute_io_wgt_rd_data_bits_1_8 = load_io_wgt_rd_data_bits_1_8; // @[Core.scala 100:18:@24704.4]
  assign compute_io_wgt_rd_data_bits_1_9 = load_io_wgt_rd_data_bits_1_9; // @[Core.scala 100:18:@24705.4]
  assign compute_io_wgt_rd_data_bits_1_10 = load_io_wgt_rd_data_bits_1_10; // @[Core.scala 100:18:@24706.4]
  assign compute_io_wgt_rd_data_bits_1_11 = load_io_wgt_rd_data_bits_1_11; // @[Core.scala 100:18:@24707.4]
  assign compute_io_wgt_rd_data_bits_1_12 = load_io_wgt_rd_data_bits_1_12; // @[Core.scala 100:18:@24708.4]
  assign compute_io_wgt_rd_data_bits_1_13 = load_io_wgt_rd_data_bits_1_13; // @[Core.scala 100:18:@24709.4]
  assign compute_io_wgt_rd_data_bits_1_14 = load_io_wgt_rd_data_bits_1_14; // @[Core.scala 100:18:@24710.4]
  assign compute_io_wgt_rd_data_bits_1_15 = load_io_wgt_rd_data_bits_1_15; // @[Core.scala 100:18:@24711.4]
  assign compute_io_wgt_rd_data_bits_2_0 = load_io_wgt_rd_data_bits_2_0; // @[Core.scala 100:18:@24712.4]
  assign compute_io_wgt_rd_data_bits_2_1 = load_io_wgt_rd_data_bits_2_1; // @[Core.scala 100:18:@24713.4]
  assign compute_io_wgt_rd_data_bits_2_2 = load_io_wgt_rd_data_bits_2_2; // @[Core.scala 100:18:@24714.4]
  assign compute_io_wgt_rd_data_bits_2_3 = load_io_wgt_rd_data_bits_2_3; // @[Core.scala 100:18:@24715.4]
  assign compute_io_wgt_rd_data_bits_2_4 = load_io_wgt_rd_data_bits_2_4; // @[Core.scala 100:18:@24716.4]
  assign compute_io_wgt_rd_data_bits_2_5 = load_io_wgt_rd_data_bits_2_5; // @[Core.scala 100:18:@24717.4]
  assign compute_io_wgt_rd_data_bits_2_6 = load_io_wgt_rd_data_bits_2_6; // @[Core.scala 100:18:@24718.4]
  assign compute_io_wgt_rd_data_bits_2_7 = load_io_wgt_rd_data_bits_2_7; // @[Core.scala 100:18:@24719.4]
  assign compute_io_wgt_rd_data_bits_2_8 = load_io_wgt_rd_data_bits_2_8; // @[Core.scala 100:18:@24720.4]
  assign compute_io_wgt_rd_data_bits_2_9 = load_io_wgt_rd_data_bits_2_9; // @[Core.scala 100:18:@24721.4]
  assign compute_io_wgt_rd_data_bits_2_10 = load_io_wgt_rd_data_bits_2_10; // @[Core.scala 100:18:@24722.4]
  assign compute_io_wgt_rd_data_bits_2_11 = load_io_wgt_rd_data_bits_2_11; // @[Core.scala 100:18:@24723.4]
  assign compute_io_wgt_rd_data_bits_2_12 = load_io_wgt_rd_data_bits_2_12; // @[Core.scala 100:18:@24724.4]
  assign compute_io_wgt_rd_data_bits_2_13 = load_io_wgt_rd_data_bits_2_13; // @[Core.scala 100:18:@24725.4]
  assign compute_io_wgt_rd_data_bits_2_14 = load_io_wgt_rd_data_bits_2_14; // @[Core.scala 100:18:@24726.4]
  assign compute_io_wgt_rd_data_bits_2_15 = load_io_wgt_rd_data_bits_2_15; // @[Core.scala 100:18:@24727.4]
  assign compute_io_wgt_rd_data_bits_3_0 = load_io_wgt_rd_data_bits_3_0; // @[Core.scala 100:18:@24728.4]
  assign compute_io_wgt_rd_data_bits_3_1 = load_io_wgt_rd_data_bits_3_1; // @[Core.scala 100:18:@24729.4]
  assign compute_io_wgt_rd_data_bits_3_2 = load_io_wgt_rd_data_bits_3_2; // @[Core.scala 100:18:@24730.4]
  assign compute_io_wgt_rd_data_bits_3_3 = load_io_wgt_rd_data_bits_3_3; // @[Core.scala 100:18:@24731.4]
  assign compute_io_wgt_rd_data_bits_3_4 = load_io_wgt_rd_data_bits_3_4; // @[Core.scala 100:18:@24732.4]
  assign compute_io_wgt_rd_data_bits_3_5 = load_io_wgt_rd_data_bits_3_5; // @[Core.scala 100:18:@24733.4]
  assign compute_io_wgt_rd_data_bits_3_6 = load_io_wgt_rd_data_bits_3_6; // @[Core.scala 100:18:@24734.4]
  assign compute_io_wgt_rd_data_bits_3_7 = load_io_wgt_rd_data_bits_3_7; // @[Core.scala 100:18:@24735.4]
  assign compute_io_wgt_rd_data_bits_3_8 = load_io_wgt_rd_data_bits_3_8; // @[Core.scala 100:18:@24736.4]
  assign compute_io_wgt_rd_data_bits_3_9 = load_io_wgt_rd_data_bits_3_9; // @[Core.scala 100:18:@24737.4]
  assign compute_io_wgt_rd_data_bits_3_10 = load_io_wgt_rd_data_bits_3_10; // @[Core.scala 100:18:@24738.4]
  assign compute_io_wgt_rd_data_bits_3_11 = load_io_wgt_rd_data_bits_3_11; // @[Core.scala 100:18:@24739.4]
  assign compute_io_wgt_rd_data_bits_3_12 = load_io_wgt_rd_data_bits_3_12; // @[Core.scala 100:18:@24740.4]
  assign compute_io_wgt_rd_data_bits_3_13 = load_io_wgt_rd_data_bits_3_13; // @[Core.scala 100:18:@24741.4]
  assign compute_io_wgt_rd_data_bits_3_14 = load_io_wgt_rd_data_bits_3_14; // @[Core.scala 100:18:@24742.4]
  assign compute_io_wgt_rd_data_bits_3_15 = load_io_wgt_rd_data_bits_3_15; // @[Core.scala 100:18:@24743.4]
  assign compute_io_wgt_rd_data_bits_4_0 = load_io_wgt_rd_data_bits_4_0; // @[Core.scala 100:18:@24744.4]
  assign compute_io_wgt_rd_data_bits_4_1 = load_io_wgt_rd_data_bits_4_1; // @[Core.scala 100:18:@24745.4]
  assign compute_io_wgt_rd_data_bits_4_2 = load_io_wgt_rd_data_bits_4_2; // @[Core.scala 100:18:@24746.4]
  assign compute_io_wgt_rd_data_bits_4_3 = load_io_wgt_rd_data_bits_4_3; // @[Core.scala 100:18:@24747.4]
  assign compute_io_wgt_rd_data_bits_4_4 = load_io_wgt_rd_data_bits_4_4; // @[Core.scala 100:18:@24748.4]
  assign compute_io_wgt_rd_data_bits_4_5 = load_io_wgt_rd_data_bits_4_5; // @[Core.scala 100:18:@24749.4]
  assign compute_io_wgt_rd_data_bits_4_6 = load_io_wgt_rd_data_bits_4_6; // @[Core.scala 100:18:@24750.4]
  assign compute_io_wgt_rd_data_bits_4_7 = load_io_wgt_rd_data_bits_4_7; // @[Core.scala 100:18:@24751.4]
  assign compute_io_wgt_rd_data_bits_4_8 = load_io_wgt_rd_data_bits_4_8; // @[Core.scala 100:18:@24752.4]
  assign compute_io_wgt_rd_data_bits_4_9 = load_io_wgt_rd_data_bits_4_9; // @[Core.scala 100:18:@24753.4]
  assign compute_io_wgt_rd_data_bits_4_10 = load_io_wgt_rd_data_bits_4_10; // @[Core.scala 100:18:@24754.4]
  assign compute_io_wgt_rd_data_bits_4_11 = load_io_wgt_rd_data_bits_4_11; // @[Core.scala 100:18:@24755.4]
  assign compute_io_wgt_rd_data_bits_4_12 = load_io_wgt_rd_data_bits_4_12; // @[Core.scala 100:18:@24756.4]
  assign compute_io_wgt_rd_data_bits_4_13 = load_io_wgt_rd_data_bits_4_13; // @[Core.scala 100:18:@24757.4]
  assign compute_io_wgt_rd_data_bits_4_14 = load_io_wgt_rd_data_bits_4_14; // @[Core.scala 100:18:@24758.4]
  assign compute_io_wgt_rd_data_bits_4_15 = load_io_wgt_rd_data_bits_4_15; // @[Core.scala 100:18:@24759.4]
  assign compute_io_wgt_rd_data_bits_5_0 = load_io_wgt_rd_data_bits_5_0; // @[Core.scala 100:18:@24760.4]
  assign compute_io_wgt_rd_data_bits_5_1 = load_io_wgt_rd_data_bits_5_1; // @[Core.scala 100:18:@24761.4]
  assign compute_io_wgt_rd_data_bits_5_2 = load_io_wgt_rd_data_bits_5_2; // @[Core.scala 100:18:@24762.4]
  assign compute_io_wgt_rd_data_bits_5_3 = load_io_wgt_rd_data_bits_5_3; // @[Core.scala 100:18:@24763.4]
  assign compute_io_wgt_rd_data_bits_5_4 = load_io_wgt_rd_data_bits_5_4; // @[Core.scala 100:18:@24764.4]
  assign compute_io_wgt_rd_data_bits_5_5 = load_io_wgt_rd_data_bits_5_5; // @[Core.scala 100:18:@24765.4]
  assign compute_io_wgt_rd_data_bits_5_6 = load_io_wgt_rd_data_bits_5_6; // @[Core.scala 100:18:@24766.4]
  assign compute_io_wgt_rd_data_bits_5_7 = load_io_wgt_rd_data_bits_5_7; // @[Core.scala 100:18:@24767.4]
  assign compute_io_wgt_rd_data_bits_5_8 = load_io_wgt_rd_data_bits_5_8; // @[Core.scala 100:18:@24768.4]
  assign compute_io_wgt_rd_data_bits_5_9 = load_io_wgt_rd_data_bits_5_9; // @[Core.scala 100:18:@24769.4]
  assign compute_io_wgt_rd_data_bits_5_10 = load_io_wgt_rd_data_bits_5_10; // @[Core.scala 100:18:@24770.4]
  assign compute_io_wgt_rd_data_bits_5_11 = load_io_wgt_rd_data_bits_5_11; // @[Core.scala 100:18:@24771.4]
  assign compute_io_wgt_rd_data_bits_5_12 = load_io_wgt_rd_data_bits_5_12; // @[Core.scala 100:18:@24772.4]
  assign compute_io_wgt_rd_data_bits_5_13 = load_io_wgt_rd_data_bits_5_13; // @[Core.scala 100:18:@24773.4]
  assign compute_io_wgt_rd_data_bits_5_14 = load_io_wgt_rd_data_bits_5_14; // @[Core.scala 100:18:@24774.4]
  assign compute_io_wgt_rd_data_bits_5_15 = load_io_wgt_rd_data_bits_5_15; // @[Core.scala 100:18:@24775.4]
  assign compute_io_wgt_rd_data_bits_6_0 = load_io_wgt_rd_data_bits_6_0; // @[Core.scala 100:18:@24776.4]
  assign compute_io_wgt_rd_data_bits_6_1 = load_io_wgt_rd_data_bits_6_1; // @[Core.scala 100:18:@24777.4]
  assign compute_io_wgt_rd_data_bits_6_2 = load_io_wgt_rd_data_bits_6_2; // @[Core.scala 100:18:@24778.4]
  assign compute_io_wgt_rd_data_bits_6_3 = load_io_wgt_rd_data_bits_6_3; // @[Core.scala 100:18:@24779.4]
  assign compute_io_wgt_rd_data_bits_6_4 = load_io_wgt_rd_data_bits_6_4; // @[Core.scala 100:18:@24780.4]
  assign compute_io_wgt_rd_data_bits_6_5 = load_io_wgt_rd_data_bits_6_5; // @[Core.scala 100:18:@24781.4]
  assign compute_io_wgt_rd_data_bits_6_6 = load_io_wgt_rd_data_bits_6_6; // @[Core.scala 100:18:@24782.4]
  assign compute_io_wgt_rd_data_bits_6_7 = load_io_wgt_rd_data_bits_6_7; // @[Core.scala 100:18:@24783.4]
  assign compute_io_wgt_rd_data_bits_6_8 = load_io_wgt_rd_data_bits_6_8; // @[Core.scala 100:18:@24784.4]
  assign compute_io_wgt_rd_data_bits_6_9 = load_io_wgt_rd_data_bits_6_9; // @[Core.scala 100:18:@24785.4]
  assign compute_io_wgt_rd_data_bits_6_10 = load_io_wgt_rd_data_bits_6_10; // @[Core.scala 100:18:@24786.4]
  assign compute_io_wgt_rd_data_bits_6_11 = load_io_wgt_rd_data_bits_6_11; // @[Core.scala 100:18:@24787.4]
  assign compute_io_wgt_rd_data_bits_6_12 = load_io_wgt_rd_data_bits_6_12; // @[Core.scala 100:18:@24788.4]
  assign compute_io_wgt_rd_data_bits_6_13 = load_io_wgt_rd_data_bits_6_13; // @[Core.scala 100:18:@24789.4]
  assign compute_io_wgt_rd_data_bits_6_14 = load_io_wgt_rd_data_bits_6_14; // @[Core.scala 100:18:@24790.4]
  assign compute_io_wgt_rd_data_bits_6_15 = load_io_wgt_rd_data_bits_6_15; // @[Core.scala 100:18:@24791.4]
  assign compute_io_wgt_rd_data_bits_7_0 = load_io_wgt_rd_data_bits_7_0; // @[Core.scala 100:18:@24792.4]
  assign compute_io_wgt_rd_data_bits_7_1 = load_io_wgt_rd_data_bits_7_1; // @[Core.scala 100:18:@24793.4]
  assign compute_io_wgt_rd_data_bits_7_2 = load_io_wgt_rd_data_bits_7_2; // @[Core.scala 100:18:@24794.4]
  assign compute_io_wgt_rd_data_bits_7_3 = load_io_wgt_rd_data_bits_7_3; // @[Core.scala 100:18:@24795.4]
  assign compute_io_wgt_rd_data_bits_7_4 = load_io_wgt_rd_data_bits_7_4; // @[Core.scala 100:18:@24796.4]
  assign compute_io_wgt_rd_data_bits_7_5 = load_io_wgt_rd_data_bits_7_5; // @[Core.scala 100:18:@24797.4]
  assign compute_io_wgt_rd_data_bits_7_6 = load_io_wgt_rd_data_bits_7_6; // @[Core.scala 100:18:@24798.4]
  assign compute_io_wgt_rd_data_bits_7_7 = load_io_wgt_rd_data_bits_7_7; // @[Core.scala 100:18:@24799.4]
  assign compute_io_wgt_rd_data_bits_7_8 = load_io_wgt_rd_data_bits_7_8; // @[Core.scala 100:18:@24800.4]
  assign compute_io_wgt_rd_data_bits_7_9 = load_io_wgt_rd_data_bits_7_9; // @[Core.scala 100:18:@24801.4]
  assign compute_io_wgt_rd_data_bits_7_10 = load_io_wgt_rd_data_bits_7_10; // @[Core.scala 100:18:@24802.4]
  assign compute_io_wgt_rd_data_bits_7_11 = load_io_wgt_rd_data_bits_7_11; // @[Core.scala 100:18:@24803.4]
  assign compute_io_wgt_rd_data_bits_7_12 = load_io_wgt_rd_data_bits_7_12; // @[Core.scala 100:18:@24804.4]
  assign compute_io_wgt_rd_data_bits_7_13 = load_io_wgt_rd_data_bits_7_13; // @[Core.scala 100:18:@24805.4]
  assign compute_io_wgt_rd_data_bits_7_14 = load_io_wgt_rd_data_bits_7_14; // @[Core.scala 100:18:@24806.4]
  assign compute_io_wgt_rd_data_bits_7_15 = load_io_wgt_rd_data_bits_7_15; // @[Core.scala 100:18:@24807.4]
  assign compute_io_wgt_rd_data_bits_8_0 = load_io_wgt_rd_data_bits_8_0; // @[Core.scala 100:18:@24808.4]
  assign compute_io_wgt_rd_data_bits_8_1 = load_io_wgt_rd_data_bits_8_1; // @[Core.scala 100:18:@24809.4]
  assign compute_io_wgt_rd_data_bits_8_2 = load_io_wgt_rd_data_bits_8_2; // @[Core.scala 100:18:@24810.4]
  assign compute_io_wgt_rd_data_bits_8_3 = load_io_wgt_rd_data_bits_8_3; // @[Core.scala 100:18:@24811.4]
  assign compute_io_wgt_rd_data_bits_8_4 = load_io_wgt_rd_data_bits_8_4; // @[Core.scala 100:18:@24812.4]
  assign compute_io_wgt_rd_data_bits_8_5 = load_io_wgt_rd_data_bits_8_5; // @[Core.scala 100:18:@24813.4]
  assign compute_io_wgt_rd_data_bits_8_6 = load_io_wgt_rd_data_bits_8_6; // @[Core.scala 100:18:@24814.4]
  assign compute_io_wgt_rd_data_bits_8_7 = load_io_wgt_rd_data_bits_8_7; // @[Core.scala 100:18:@24815.4]
  assign compute_io_wgt_rd_data_bits_8_8 = load_io_wgt_rd_data_bits_8_8; // @[Core.scala 100:18:@24816.4]
  assign compute_io_wgt_rd_data_bits_8_9 = load_io_wgt_rd_data_bits_8_9; // @[Core.scala 100:18:@24817.4]
  assign compute_io_wgt_rd_data_bits_8_10 = load_io_wgt_rd_data_bits_8_10; // @[Core.scala 100:18:@24818.4]
  assign compute_io_wgt_rd_data_bits_8_11 = load_io_wgt_rd_data_bits_8_11; // @[Core.scala 100:18:@24819.4]
  assign compute_io_wgt_rd_data_bits_8_12 = load_io_wgt_rd_data_bits_8_12; // @[Core.scala 100:18:@24820.4]
  assign compute_io_wgt_rd_data_bits_8_13 = load_io_wgt_rd_data_bits_8_13; // @[Core.scala 100:18:@24821.4]
  assign compute_io_wgt_rd_data_bits_8_14 = load_io_wgt_rd_data_bits_8_14; // @[Core.scala 100:18:@24822.4]
  assign compute_io_wgt_rd_data_bits_8_15 = load_io_wgt_rd_data_bits_8_15; // @[Core.scala 100:18:@24823.4]
  assign compute_io_wgt_rd_data_bits_9_0 = load_io_wgt_rd_data_bits_9_0; // @[Core.scala 100:18:@24824.4]
  assign compute_io_wgt_rd_data_bits_9_1 = load_io_wgt_rd_data_bits_9_1; // @[Core.scala 100:18:@24825.4]
  assign compute_io_wgt_rd_data_bits_9_2 = load_io_wgt_rd_data_bits_9_2; // @[Core.scala 100:18:@24826.4]
  assign compute_io_wgt_rd_data_bits_9_3 = load_io_wgt_rd_data_bits_9_3; // @[Core.scala 100:18:@24827.4]
  assign compute_io_wgt_rd_data_bits_9_4 = load_io_wgt_rd_data_bits_9_4; // @[Core.scala 100:18:@24828.4]
  assign compute_io_wgt_rd_data_bits_9_5 = load_io_wgt_rd_data_bits_9_5; // @[Core.scala 100:18:@24829.4]
  assign compute_io_wgt_rd_data_bits_9_6 = load_io_wgt_rd_data_bits_9_6; // @[Core.scala 100:18:@24830.4]
  assign compute_io_wgt_rd_data_bits_9_7 = load_io_wgt_rd_data_bits_9_7; // @[Core.scala 100:18:@24831.4]
  assign compute_io_wgt_rd_data_bits_9_8 = load_io_wgt_rd_data_bits_9_8; // @[Core.scala 100:18:@24832.4]
  assign compute_io_wgt_rd_data_bits_9_9 = load_io_wgt_rd_data_bits_9_9; // @[Core.scala 100:18:@24833.4]
  assign compute_io_wgt_rd_data_bits_9_10 = load_io_wgt_rd_data_bits_9_10; // @[Core.scala 100:18:@24834.4]
  assign compute_io_wgt_rd_data_bits_9_11 = load_io_wgt_rd_data_bits_9_11; // @[Core.scala 100:18:@24835.4]
  assign compute_io_wgt_rd_data_bits_9_12 = load_io_wgt_rd_data_bits_9_12; // @[Core.scala 100:18:@24836.4]
  assign compute_io_wgt_rd_data_bits_9_13 = load_io_wgt_rd_data_bits_9_13; // @[Core.scala 100:18:@24837.4]
  assign compute_io_wgt_rd_data_bits_9_14 = load_io_wgt_rd_data_bits_9_14; // @[Core.scala 100:18:@24838.4]
  assign compute_io_wgt_rd_data_bits_9_15 = load_io_wgt_rd_data_bits_9_15; // @[Core.scala 100:18:@24839.4]
  assign compute_io_wgt_rd_data_bits_10_0 = load_io_wgt_rd_data_bits_10_0; // @[Core.scala 100:18:@24840.4]
  assign compute_io_wgt_rd_data_bits_10_1 = load_io_wgt_rd_data_bits_10_1; // @[Core.scala 100:18:@24841.4]
  assign compute_io_wgt_rd_data_bits_10_2 = load_io_wgt_rd_data_bits_10_2; // @[Core.scala 100:18:@24842.4]
  assign compute_io_wgt_rd_data_bits_10_3 = load_io_wgt_rd_data_bits_10_3; // @[Core.scala 100:18:@24843.4]
  assign compute_io_wgt_rd_data_bits_10_4 = load_io_wgt_rd_data_bits_10_4; // @[Core.scala 100:18:@24844.4]
  assign compute_io_wgt_rd_data_bits_10_5 = load_io_wgt_rd_data_bits_10_5; // @[Core.scala 100:18:@24845.4]
  assign compute_io_wgt_rd_data_bits_10_6 = load_io_wgt_rd_data_bits_10_6; // @[Core.scala 100:18:@24846.4]
  assign compute_io_wgt_rd_data_bits_10_7 = load_io_wgt_rd_data_bits_10_7; // @[Core.scala 100:18:@24847.4]
  assign compute_io_wgt_rd_data_bits_10_8 = load_io_wgt_rd_data_bits_10_8; // @[Core.scala 100:18:@24848.4]
  assign compute_io_wgt_rd_data_bits_10_9 = load_io_wgt_rd_data_bits_10_9; // @[Core.scala 100:18:@24849.4]
  assign compute_io_wgt_rd_data_bits_10_10 = load_io_wgt_rd_data_bits_10_10; // @[Core.scala 100:18:@24850.4]
  assign compute_io_wgt_rd_data_bits_10_11 = load_io_wgt_rd_data_bits_10_11; // @[Core.scala 100:18:@24851.4]
  assign compute_io_wgt_rd_data_bits_10_12 = load_io_wgt_rd_data_bits_10_12; // @[Core.scala 100:18:@24852.4]
  assign compute_io_wgt_rd_data_bits_10_13 = load_io_wgt_rd_data_bits_10_13; // @[Core.scala 100:18:@24853.4]
  assign compute_io_wgt_rd_data_bits_10_14 = load_io_wgt_rd_data_bits_10_14; // @[Core.scala 100:18:@24854.4]
  assign compute_io_wgt_rd_data_bits_10_15 = load_io_wgt_rd_data_bits_10_15; // @[Core.scala 100:18:@24855.4]
  assign compute_io_wgt_rd_data_bits_11_0 = load_io_wgt_rd_data_bits_11_0; // @[Core.scala 100:18:@24856.4]
  assign compute_io_wgt_rd_data_bits_11_1 = load_io_wgt_rd_data_bits_11_1; // @[Core.scala 100:18:@24857.4]
  assign compute_io_wgt_rd_data_bits_11_2 = load_io_wgt_rd_data_bits_11_2; // @[Core.scala 100:18:@24858.4]
  assign compute_io_wgt_rd_data_bits_11_3 = load_io_wgt_rd_data_bits_11_3; // @[Core.scala 100:18:@24859.4]
  assign compute_io_wgt_rd_data_bits_11_4 = load_io_wgt_rd_data_bits_11_4; // @[Core.scala 100:18:@24860.4]
  assign compute_io_wgt_rd_data_bits_11_5 = load_io_wgt_rd_data_bits_11_5; // @[Core.scala 100:18:@24861.4]
  assign compute_io_wgt_rd_data_bits_11_6 = load_io_wgt_rd_data_bits_11_6; // @[Core.scala 100:18:@24862.4]
  assign compute_io_wgt_rd_data_bits_11_7 = load_io_wgt_rd_data_bits_11_7; // @[Core.scala 100:18:@24863.4]
  assign compute_io_wgt_rd_data_bits_11_8 = load_io_wgt_rd_data_bits_11_8; // @[Core.scala 100:18:@24864.4]
  assign compute_io_wgt_rd_data_bits_11_9 = load_io_wgt_rd_data_bits_11_9; // @[Core.scala 100:18:@24865.4]
  assign compute_io_wgt_rd_data_bits_11_10 = load_io_wgt_rd_data_bits_11_10; // @[Core.scala 100:18:@24866.4]
  assign compute_io_wgt_rd_data_bits_11_11 = load_io_wgt_rd_data_bits_11_11; // @[Core.scala 100:18:@24867.4]
  assign compute_io_wgt_rd_data_bits_11_12 = load_io_wgt_rd_data_bits_11_12; // @[Core.scala 100:18:@24868.4]
  assign compute_io_wgt_rd_data_bits_11_13 = load_io_wgt_rd_data_bits_11_13; // @[Core.scala 100:18:@24869.4]
  assign compute_io_wgt_rd_data_bits_11_14 = load_io_wgt_rd_data_bits_11_14; // @[Core.scala 100:18:@24870.4]
  assign compute_io_wgt_rd_data_bits_11_15 = load_io_wgt_rd_data_bits_11_15; // @[Core.scala 100:18:@24871.4]
  assign compute_io_wgt_rd_data_bits_12_0 = load_io_wgt_rd_data_bits_12_0; // @[Core.scala 100:18:@24872.4]
  assign compute_io_wgt_rd_data_bits_12_1 = load_io_wgt_rd_data_bits_12_1; // @[Core.scala 100:18:@24873.4]
  assign compute_io_wgt_rd_data_bits_12_2 = load_io_wgt_rd_data_bits_12_2; // @[Core.scala 100:18:@24874.4]
  assign compute_io_wgt_rd_data_bits_12_3 = load_io_wgt_rd_data_bits_12_3; // @[Core.scala 100:18:@24875.4]
  assign compute_io_wgt_rd_data_bits_12_4 = load_io_wgt_rd_data_bits_12_4; // @[Core.scala 100:18:@24876.4]
  assign compute_io_wgt_rd_data_bits_12_5 = load_io_wgt_rd_data_bits_12_5; // @[Core.scala 100:18:@24877.4]
  assign compute_io_wgt_rd_data_bits_12_6 = load_io_wgt_rd_data_bits_12_6; // @[Core.scala 100:18:@24878.4]
  assign compute_io_wgt_rd_data_bits_12_7 = load_io_wgt_rd_data_bits_12_7; // @[Core.scala 100:18:@24879.4]
  assign compute_io_wgt_rd_data_bits_12_8 = load_io_wgt_rd_data_bits_12_8; // @[Core.scala 100:18:@24880.4]
  assign compute_io_wgt_rd_data_bits_12_9 = load_io_wgt_rd_data_bits_12_9; // @[Core.scala 100:18:@24881.4]
  assign compute_io_wgt_rd_data_bits_12_10 = load_io_wgt_rd_data_bits_12_10; // @[Core.scala 100:18:@24882.4]
  assign compute_io_wgt_rd_data_bits_12_11 = load_io_wgt_rd_data_bits_12_11; // @[Core.scala 100:18:@24883.4]
  assign compute_io_wgt_rd_data_bits_12_12 = load_io_wgt_rd_data_bits_12_12; // @[Core.scala 100:18:@24884.4]
  assign compute_io_wgt_rd_data_bits_12_13 = load_io_wgt_rd_data_bits_12_13; // @[Core.scala 100:18:@24885.4]
  assign compute_io_wgt_rd_data_bits_12_14 = load_io_wgt_rd_data_bits_12_14; // @[Core.scala 100:18:@24886.4]
  assign compute_io_wgt_rd_data_bits_12_15 = load_io_wgt_rd_data_bits_12_15; // @[Core.scala 100:18:@24887.4]
  assign compute_io_wgt_rd_data_bits_13_0 = load_io_wgt_rd_data_bits_13_0; // @[Core.scala 100:18:@24888.4]
  assign compute_io_wgt_rd_data_bits_13_1 = load_io_wgt_rd_data_bits_13_1; // @[Core.scala 100:18:@24889.4]
  assign compute_io_wgt_rd_data_bits_13_2 = load_io_wgt_rd_data_bits_13_2; // @[Core.scala 100:18:@24890.4]
  assign compute_io_wgt_rd_data_bits_13_3 = load_io_wgt_rd_data_bits_13_3; // @[Core.scala 100:18:@24891.4]
  assign compute_io_wgt_rd_data_bits_13_4 = load_io_wgt_rd_data_bits_13_4; // @[Core.scala 100:18:@24892.4]
  assign compute_io_wgt_rd_data_bits_13_5 = load_io_wgt_rd_data_bits_13_5; // @[Core.scala 100:18:@24893.4]
  assign compute_io_wgt_rd_data_bits_13_6 = load_io_wgt_rd_data_bits_13_6; // @[Core.scala 100:18:@24894.4]
  assign compute_io_wgt_rd_data_bits_13_7 = load_io_wgt_rd_data_bits_13_7; // @[Core.scala 100:18:@24895.4]
  assign compute_io_wgt_rd_data_bits_13_8 = load_io_wgt_rd_data_bits_13_8; // @[Core.scala 100:18:@24896.4]
  assign compute_io_wgt_rd_data_bits_13_9 = load_io_wgt_rd_data_bits_13_9; // @[Core.scala 100:18:@24897.4]
  assign compute_io_wgt_rd_data_bits_13_10 = load_io_wgt_rd_data_bits_13_10; // @[Core.scala 100:18:@24898.4]
  assign compute_io_wgt_rd_data_bits_13_11 = load_io_wgt_rd_data_bits_13_11; // @[Core.scala 100:18:@24899.4]
  assign compute_io_wgt_rd_data_bits_13_12 = load_io_wgt_rd_data_bits_13_12; // @[Core.scala 100:18:@24900.4]
  assign compute_io_wgt_rd_data_bits_13_13 = load_io_wgt_rd_data_bits_13_13; // @[Core.scala 100:18:@24901.4]
  assign compute_io_wgt_rd_data_bits_13_14 = load_io_wgt_rd_data_bits_13_14; // @[Core.scala 100:18:@24902.4]
  assign compute_io_wgt_rd_data_bits_13_15 = load_io_wgt_rd_data_bits_13_15; // @[Core.scala 100:18:@24903.4]
  assign compute_io_wgt_rd_data_bits_14_0 = load_io_wgt_rd_data_bits_14_0; // @[Core.scala 100:18:@24904.4]
  assign compute_io_wgt_rd_data_bits_14_1 = load_io_wgt_rd_data_bits_14_1; // @[Core.scala 100:18:@24905.4]
  assign compute_io_wgt_rd_data_bits_14_2 = load_io_wgt_rd_data_bits_14_2; // @[Core.scala 100:18:@24906.4]
  assign compute_io_wgt_rd_data_bits_14_3 = load_io_wgt_rd_data_bits_14_3; // @[Core.scala 100:18:@24907.4]
  assign compute_io_wgt_rd_data_bits_14_4 = load_io_wgt_rd_data_bits_14_4; // @[Core.scala 100:18:@24908.4]
  assign compute_io_wgt_rd_data_bits_14_5 = load_io_wgt_rd_data_bits_14_5; // @[Core.scala 100:18:@24909.4]
  assign compute_io_wgt_rd_data_bits_14_6 = load_io_wgt_rd_data_bits_14_6; // @[Core.scala 100:18:@24910.4]
  assign compute_io_wgt_rd_data_bits_14_7 = load_io_wgt_rd_data_bits_14_7; // @[Core.scala 100:18:@24911.4]
  assign compute_io_wgt_rd_data_bits_14_8 = load_io_wgt_rd_data_bits_14_8; // @[Core.scala 100:18:@24912.4]
  assign compute_io_wgt_rd_data_bits_14_9 = load_io_wgt_rd_data_bits_14_9; // @[Core.scala 100:18:@24913.4]
  assign compute_io_wgt_rd_data_bits_14_10 = load_io_wgt_rd_data_bits_14_10; // @[Core.scala 100:18:@24914.4]
  assign compute_io_wgt_rd_data_bits_14_11 = load_io_wgt_rd_data_bits_14_11; // @[Core.scala 100:18:@24915.4]
  assign compute_io_wgt_rd_data_bits_14_12 = load_io_wgt_rd_data_bits_14_12; // @[Core.scala 100:18:@24916.4]
  assign compute_io_wgt_rd_data_bits_14_13 = load_io_wgt_rd_data_bits_14_13; // @[Core.scala 100:18:@24917.4]
  assign compute_io_wgt_rd_data_bits_14_14 = load_io_wgt_rd_data_bits_14_14; // @[Core.scala 100:18:@24918.4]
  assign compute_io_wgt_rd_data_bits_14_15 = load_io_wgt_rd_data_bits_14_15; // @[Core.scala 100:18:@24919.4]
  assign compute_io_wgt_rd_data_bits_15_0 = load_io_wgt_rd_data_bits_15_0; // @[Core.scala 100:18:@24920.4]
  assign compute_io_wgt_rd_data_bits_15_1 = load_io_wgt_rd_data_bits_15_1; // @[Core.scala 100:18:@24921.4]
  assign compute_io_wgt_rd_data_bits_15_2 = load_io_wgt_rd_data_bits_15_2; // @[Core.scala 100:18:@24922.4]
  assign compute_io_wgt_rd_data_bits_15_3 = load_io_wgt_rd_data_bits_15_3; // @[Core.scala 100:18:@24923.4]
  assign compute_io_wgt_rd_data_bits_15_4 = load_io_wgt_rd_data_bits_15_4; // @[Core.scala 100:18:@24924.4]
  assign compute_io_wgt_rd_data_bits_15_5 = load_io_wgt_rd_data_bits_15_5; // @[Core.scala 100:18:@24925.4]
  assign compute_io_wgt_rd_data_bits_15_6 = load_io_wgt_rd_data_bits_15_6; // @[Core.scala 100:18:@24926.4]
  assign compute_io_wgt_rd_data_bits_15_7 = load_io_wgt_rd_data_bits_15_7; // @[Core.scala 100:18:@24927.4]
  assign compute_io_wgt_rd_data_bits_15_8 = load_io_wgt_rd_data_bits_15_8; // @[Core.scala 100:18:@24928.4]
  assign compute_io_wgt_rd_data_bits_15_9 = load_io_wgt_rd_data_bits_15_9; // @[Core.scala 100:18:@24929.4]
  assign compute_io_wgt_rd_data_bits_15_10 = load_io_wgt_rd_data_bits_15_10; // @[Core.scala 100:18:@24930.4]
  assign compute_io_wgt_rd_data_bits_15_11 = load_io_wgt_rd_data_bits_15_11; // @[Core.scala 100:18:@24931.4]
  assign compute_io_wgt_rd_data_bits_15_12 = load_io_wgt_rd_data_bits_15_12; // @[Core.scala 100:18:@24932.4]
  assign compute_io_wgt_rd_data_bits_15_13 = load_io_wgt_rd_data_bits_15_13; // @[Core.scala 100:18:@24933.4]
  assign compute_io_wgt_rd_data_bits_15_14 = load_io_wgt_rd_data_bits_15_14; // @[Core.scala 100:18:@24934.4]
  assign compute_io_wgt_rd_data_bits_15_15 = load_io_wgt_rd_data_bits_15_15; // @[Core.scala 100:18:@24935.4]
  assign store_clock = clock; // @[:@24321.4]
  assign store_reset = reset; // @[:@24322.4]
  assign store_io_i_post = compute_io_o_post_1; // @[Core.scala 105:19:@24939.4]
  assign store_io_inst_valid = fetch_io_inst_st_valid; // @[Core.scala 106:17:@24941.4]
  assign store_io_inst_bits = fetch_io_inst_st_bits; // @[Core.scala 106:17:@24940.4]
  assign store_io_out_baddr = io_vcr_ptrs_5; // @[Core.scala 107:22:@24943.4]
  assign store_io_vme_wr_cmd_ready = io_vme_wr_0_cmd_ready; // @[Core.scala 78:16:@24368.4]
  assign store_io_vme_wr_data_ready = io_vme_wr_0_data_ready; // @[Core.scala 78:16:@24364.4]
  assign store_io_vme_wr_ack = io_vme_wr_0_ack; // @[Core.scala 78:16:@24361.4]
  assign store_io_out_wr_valid = compute_io_out_wr_valid; // @[Core.scala 108:16:@24961.4]
  assign store_io_out_wr_bits_idx = compute_io_out_wr_bits_idx; // @[Core.scala 108:16:@24960.4]
  assign store_io_out_wr_bits_data_0_0 = compute_io_out_wr_bits_data_0_0; // @[Core.scala 108:16:@24944.4]
  assign store_io_out_wr_bits_data_0_1 = compute_io_out_wr_bits_data_0_1; // @[Core.scala 108:16:@24945.4]
  assign store_io_out_wr_bits_data_0_2 = compute_io_out_wr_bits_data_0_2; // @[Core.scala 108:16:@24946.4]
  assign store_io_out_wr_bits_data_0_3 = compute_io_out_wr_bits_data_0_3; // @[Core.scala 108:16:@24947.4]
  assign store_io_out_wr_bits_data_0_4 = compute_io_out_wr_bits_data_0_4; // @[Core.scala 108:16:@24948.4]
  assign store_io_out_wr_bits_data_0_5 = compute_io_out_wr_bits_data_0_5; // @[Core.scala 108:16:@24949.4]
  assign store_io_out_wr_bits_data_0_6 = compute_io_out_wr_bits_data_0_6; // @[Core.scala 108:16:@24950.4]
  assign store_io_out_wr_bits_data_0_7 = compute_io_out_wr_bits_data_0_7; // @[Core.scala 108:16:@24951.4]
  assign store_io_out_wr_bits_data_0_8 = compute_io_out_wr_bits_data_0_8; // @[Core.scala 108:16:@24952.4]
  assign store_io_out_wr_bits_data_0_9 = compute_io_out_wr_bits_data_0_9; // @[Core.scala 108:16:@24953.4]
  assign store_io_out_wr_bits_data_0_10 = compute_io_out_wr_bits_data_0_10; // @[Core.scala 108:16:@24954.4]
  assign store_io_out_wr_bits_data_0_11 = compute_io_out_wr_bits_data_0_11; // @[Core.scala 108:16:@24955.4]
  assign store_io_out_wr_bits_data_0_12 = compute_io_out_wr_bits_data_0_12; // @[Core.scala 108:16:@24956.4]
  assign store_io_out_wr_bits_data_0_13 = compute_io_out_wr_bits_data_0_13; // @[Core.scala 108:16:@24957.4]
  assign store_io_out_wr_bits_data_0_14 = compute_io_out_wr_bits_data_0_14; // @[Core.scala 108:16:@24958.4]
  assign store_io_out_wr_bits_data_0_15 = compute_io_out_wr_bits_data_0_15; // @[Core.scala 108:16:@24959.4]
  assign ecounters_clock = clock; // @[:@24324.4]
  assign ecounters_reset = reset; // @[:@24325.4]
  assign ecounters_io_launch = io_vcr_launch; // @[Core.scala 111:23:@24981.4]
  assign ecounters_io_finish = compute_io_finish; // @[Core.scala 112:23:@24982.4]
  assign ecounters_io_acc_wr_event = compute_io_acc_wr_event; // @[Core.scala 115:29:@24987.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  finish = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    finish <= compute_io_finish;
  end
endmodule
module VTAShell( // @[:@24992.2]
  input         clock, // @[:@24993.4]
  input         reset, // @[:@24994.4]
  output        io_host_aw_ready, // @[:@24995.4]
  input         io_host_aw_valid, // @[:@24995.4]
  input  [15:0] io_host_aw_bits_addr, // @[:@24995.4]
  output        io_host_w_ready, // @[:@24995.4]
  input         io_host_w_valid, // @[:@24995.4]
  input  [31:0] io_host_w_bits_data, // @[:@24995.4]
  input         io_host_b_ready, // @[:@24995.4]
  output        io_host_b_valid, // @[:@24995.4]
  output        io_host_ar_ready, // @[:@24995.4]
  input         io_host_ar_valid, // @[:@24995.4]
  input  [15:0] io_host_ar_bits_addr, // @[:@24995.4]
  input         io_host_r_ready, // @[:@24995.4]
  output        io_host_r_valid, // @[:@24995.4]
  output [31:0] io_host_r_bits_data, // @[:@24995.4]
  input         io_mem_aw_ready, // @[:@24995.4]
  output        io_mem_aw_valid, // @[:@24995.4]
  output [31:0] io_mem_aw_bits_addr, // @[:@24995.4]
  output [7:0]  io_mem_aw_bits_len, // @[:@24995.4]
  input         io_mem_w_ready, // @[:@24995.4]
  output        io_mem_w_valid, // @[:@24995.4]
  output [63:0] io_mem_w_bits_data, // @[:@24995.4]
  output        io_mem_w_bits_last, // @[:@24995.4]
  input         io_mem_b_valid, // @[:@24995.4]
  input         io_mem_ar_ready, // @[:@24995.4]
  output        io_mem_ar_valid, // @[:@24995.4]
  output [31:0] io_mem_ar_bits_addr, // @[:@24995.4]
  output [7:0]  io_mem_ar_bits_len, // @[:@24995.4]
  output        io_mem_r_ready, // @[:@24995.4]
  input         io_mem_r_valid, // @[:@24995.4]
  input  [63:0] io_mem_r_bits_data, // @[:@24995.4]
  input         io_mem_r_bits_last // @[:@24995.4]
);
  wire  vcr_clock; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_reset; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_aw_ready; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_aw_valid; // @[VTAShell.scala 48:19:@24997.4]
  wire [15:0] vcr_io_host_aw_bits_addr; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_w_ready; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_w_valid; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_host_w_bits_data; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_b_ready; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_b_valid; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_ar_ready; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_ar_valid; // @[VTAShell.scala 48:19:@24997.4]
  wire [15:0] vcr_io_host_ar_bits_addr; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_r_ready; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_host_r_valid; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_host_r_bits_data; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_vcr_launch; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_vcr_finish; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_vcr_ecnt_0_valid; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_vcr_ecnt_0_bits; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_vcr_vals_0; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_vcr_ptrs_0; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_vcr_ptrs_1; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_vcr_ptrs_2; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_vcr_ptrs_3; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_vcr_ptrs_4; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_vcr_ptrs_5; // @[VTAShell.scala 48:19:@24997.4]
  wire  vcr_io_vcr_ucnt_0_valid; // @[VTAShell.scala 48:19:@24997.4]
  wire [31:0] vcr_io_vcr_ucnt_0_bits; // @[VTAShell.scala 48:19:@24997.4]
  wire  vme_clock; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_reset; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_aw_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_aw_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [31:0] vme_io_mem_aw_bits_addr; // @[VTAShell.scala 49:19:@25000.4]
  wire [7:0] vme_io_mem_aw_bits_len; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_w_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_w_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [63:0] vme_io_mem_w_bits_data; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_w_bits_last; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_b_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_b_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_ar_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_ar_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [31:0] vme_io_mem_ar_bits_addr; // @[VTAShell.scala 49:19:@25000.4]
  wire [7:0] vme_io_mem_ar_bits_len; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_r_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_r_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [63:0] vme_io_mem_r_bits_data; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_mem_r_bits_last; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_0_cmd_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_0_cmd_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [31:0] vme_io_vme_rd_0_cmd_bits_addr; // @[VTAShell.scala 49:19:@25000.4]
  wire [7:0] vme_io_vme_rd_0_cmd_bits_len; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_0_data_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_0_data_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [63:0] vme_io_vme_rd_0_data_bits; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_1_cmd_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_1_cmd_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [31:0] vme_io_vme_rd_1_cmd_bits_addr; // @[VTAShell.scala 49:19:@25000.4]
  wire [7:0] vme_io_vme_rd_1_cmd_bits_len; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_1_data_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_1_data_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [63:0] vme_io_vme_rd_1_data_bits; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_2_cmd_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_2_cmd_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [31:0] vme_io_vme_rd_2_cmd_bits_addr; // @[VTAShell.scala 49:19:@25000.4]
  wire [7:0] vme_io_vme_rd_2_cmd_bits_len; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_2_data_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_2_data_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [63:0] vme_io_vme_rd_2_data_bits; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_3_cmd_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_3_cmd_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [31:0] vme_io_vme_rd_3_cmd_bits_addr; // @[VTAShell.scala 49:19:@25000.4]
  wire [7:0] vme_io_vme_rd_3_cmd_bits_len; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_3_data_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_3_data_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [63:0] vme_io_vme_rd_3_data_bits; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_4_cmd_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_4_cmd_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [31:0] vme_io_vme_rd_4_cmd_bits_addr; // @[VTAShell.scala 49:19:@25000.4]
  wire [7:0] vme_io_vme_rd_4_cmd_bits_len; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_4_data_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_rd_4_data_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [63:0] vme_io_vme_rd_4_data_bits; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_wr_0_cmd_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_wr_0_cmd_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [31:0] vme_io_vme_wr_0_cmd_bits_addr; // @[VTAShell.scala 49:19:@25000.4]
  wire [7:0] vme_io_vme_wr_0_cmd_bits_len; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_wr_0_data_ready; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_wr_0_data_valid; // @[VTAShell.scala 49:19:@25000.4]
  wire [63:0] vme_io_vme_wr_0_data_bits; // @[VTAShell.scala 49:19:@25000.4]
  wire  vme_io_vme_wr_0_ack; // @[VTAShell.scala 49:19:@25000.4]
  wire  core_clock; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_reset; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vcr_launch; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vcr_finish; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vcr_ecnt_0_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vcr_ecnt_0_bits; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vcr_vals_0; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vcr_ptrs_0; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vcr_ptrs_1; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vcr_ptrs_2; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vcr_ptrs_3; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vcr_ptrs_4; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vcr_ptrs_5; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vcr_ucnt_0_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vcr_ucnt_0_bits; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_0_cmd_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_0_cmd_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vme_rd_0_cmd_bits_addr; // @[VTAShell.scala 50:20:@25003.4]
  wire [7:0] core_io_vme_rd_0_cmd_bits_len; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_0_data_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_0_data_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [63:0] core_io_vme_rd_0_data_bits; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_1_cmd_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_1_cmd_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vme_rd_1_cmd_bits_addr; // @[VTAShell.scala 50:20:@25003.4]
  wire [7:0] core_io_vme_rd_1_cmd_bits_len; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_1_data_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_1_data_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [63:0] core_io_vme_rd_1_data_bits; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_2_cmd_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_2_cmd_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vme_rd_2_cmd_bits_addr; // @[VTAShell.scala 50:20:@25003.4]
  wire [7:0] core_io_vme_rd_2_cmd_bits_len; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_2_data_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_2_data_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [63:0] core_io_vme_rd_2_data_bits; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_3_cmd_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_3_cmd_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vme_rd_3_cmd_bits_addr; // @[VTAShell.scala 50:20:@25003.4]
  wire [7:0] core_io_vme_rd_3_cmd_bits_len; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_3_data_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_3_data_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [63:0] core_io_vme_rd_3_data_bits; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_4_cmd_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_4_cmd_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vme_rd_4_cmd_bits_addr; // @[VTAShell.scala 50:20:@25003.4]
  wire [7:0] core_io_vme_rd_4_cmd_bits_len; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_4_data_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_rd_4_data_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [63:0] core_io_vme_rd_4_data_bits; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_wr_0_cmd_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_wr_0_cmd_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [31:0] core_io_vme_wr_0_cmd_bits_addr; // @[VTAShell.scala 50:20:@25003.4]
  wire [7:0] core_io_vme_wr_0_cmd_bits_len; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_wr_0_data_ready; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_wr_0_data_valid; // @[VTAShell.scala 50:20:@25003.4]
  wire [63:0] core_io_vme_wr_0_data_bits; // @[VTAShell.scala 50:20:@25003.4]
  wire  core_io_vme_wr_0_ack; // @[VTAShell.scala 50:20:@25003.4]
  VCR vcr ( // @[VTAShell.scala 48:19:@24997.4]
    .clock(vcr_clock),
    .reset(vcr_reset),
    .io_host_aw_ready(vcr_io_host_aw_ready),
    .io_host_aw_valid(vcr_io_host_aw_valid),
    .io_host_aw_bits_addr(vcr_io_host_aw_bits_addr),
    .io_host_w_ready(vcr_io_host_w_ready),
    .io_host_w_valid(vcr_io_host_w_valid),
    .io_host_w_bits_data(vcr_io_host_w_bits_data),
    .io_host_b_ready(vcr_io_host_b_ready),
    .io_host_b_valid(vcr_io_host_b_valid),
    .io_host_ar_ready(vcr_io_host_ar_ready),
    .io_host_ar_valid(vcr_io_host_ar_valid),
    .io_host_ar_bits_addr(vcr_io_host_ar_bits_addr),
    .io_host_r_ready(vcr_io_host_r_ready),
    .io_host_r_valid(vcr_io_host_r_valid),
    .io_host_r_bits_data(vcr_io_host_r_bits_data),
    .io_vcr_launch(vcr_io_vcr_launch),
    .io_vcr_finish(vcr_io_vcr_finish),
    .io_vcr_ecnt_0_valid(vcr_io_vcr_ecnt_0_valid),
    .io_vcr_ecnt_0_bits(vcr_io_vcr_ecnt_0_bits),
    .io_vcr_vals_0(vcr_io_vcr_vals_0),
    .io_vcr_ptrs_0(vcr_io_vcr_ptrs_0),
    .io_vcr_ptrs_1(vcr_io_vcr_ptrs_1),
    .io_vcr_ptrs_2(vcr_io_vcr_ptrs_2),
    .io_vcr_ptrs_3(vcr_io_vcr_ptrs_3),
    .io_vcr_ptrs_4(vcr_io_vcr_ptrs_4),
    .io_vcr_ptrs_5(vcr_io_vcr_ptrs_5),
    .io_vcr_ucnt_0_valid(vcr_io_vcr_ucnt_0_valid),
    .io_vcr_ucnt_0_bits(vcr_io_vcr_ucnt_0_bits)
  );
  VME vme ( // @[VTAShell.scala 49:19:@25000.4]
    .clock(vme_clock),
    .reset(vme_reset),
    .io_mem_aw_ready(vme_io_mem_aw_ready),
    .io_mem_aw_valid(vme_io_mem_aw_valid),
    .io_mem_aw_bits_addr(vme_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(vme_io_mem_aw_bits_len),
    .io_mem_w_ready(vme_io_mem_w_ready),
    .io_mem_w_valid(vme_io_mem_w_valid),
    .io_mem_w_bits_data(vme_io_mem_w_bits_data),
    .io_mem_w_bits_last(vme_io_mem_w_bits_last),
    .io_mem_b_ready(vme_io_mem_b_ready),
    .io_mem_b_valid(vme_io_mem_b_valid),
    .io_mem_ar_ready(vme_io_mem_ar_ready),
    .io_mem_ar_valid(vme_io_mem_ar_valid),
    .io_mem_ar_bits_addr(vme_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(vme_io_mem_ar_bits_len),
    .io_mem_r_ready(vme_io_mem_r_ready),
    .io_mem_r_valid(vme_io_mem_r_valid),
    .io_mem_r_bits_data(vme_io_mem_r_bits_data),
    .io_mem_r_bits_last(vme_io_mem_r_bits_last),
    .io_vme_rd_0_cmd_ready(vme_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(vme_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(vme_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(vme_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(vme_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(vme_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits(vme_io_vme_rd_0_data_bits),
    .io_vme_rd_1_cmd_ready(vme_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(vme_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(vme_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(vme_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_data_ready(vme_io_vme_rd_1_data_ready),
    .io_vme_rd_1_data_valid(vme_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits(vme_io_vme_rd_1_data_bits),
    .io_vme_rd_2_cmd_ready(vme_io_vme_rd_2_cmd_ready),
    .io_vme_rd_2_cmd_valid(vme_io_vme_rd_2_cmd_valid),
    .io_vme_rd_2_cmd_bits_addr(vme_io_vme_rd_2_cmd_bits_addr),
    .io_vme_rd_2_cmd_bits_len(vme_io_vme_rd_2_cmd_bits_len),
    .io_vme_rd_2_data_ready(vme_io_vme_rd_2_data_ready),
    .io_vme_rd_2_data_valid(vme_io_vme_rd_2_data_valid),
    .io_vme_rd_2_data_bits(vme_io_vme_rd_2_data_bits),
    .io_vme_rd_3_cmd_ready(vme_io_vme_rd_3_cmd_ready),
    .io_vme_rd_3_cmd_valid(vme_io_vme_rd_3_cmd_valid),
    .io_vme_rd_3_cmd_bits_addr(vme_io_vme_rd_3_cmd_bits_addr),
    .io_vme_rd_3_cmd_bits_len(vme_io_vme_rd_3_cmd_bits_len),
    .io_vme_rd_3_data_ready(vme_io_vme_rd_3_data_ready),
    .io_vme_rd_3_data_valid(vme_io_vme_rd_3_data_valid),
    .io_vme_rd_3_data_bits(vme_io_vme_rd_3_data_bits),
    .io_vme_rd_4_cmd_ready(vme_io_vme_rd_4_cmd_ready),
    .io_vme_rd_4_cmd_valid(vme_io_vme_rd_4_cmd_valid),
    .io_vme_rd_4_cmd_bits_addr(vme_io_vme_rd_4_cmd_bits_addr),
    .io_vme_rd_4_cmd_bits_len(vme_io_vme_rd_4_cmd_bits_len),
    .io_vme_rd_4_data_ready(vme_io_vme_rd_4_data_ready),
    .io_vme_rd_4_data_valid(vme_io_vme_rd_4_data_valid),
    .io_vme_rd_4_data_bits(vme_io_vme_rd_4_data_bits),
    .io_vme_wr_0_cmd_ready(vme_io_vme_wr_0_cmd_ready),
    .io_vme_wr_0_cmd_valid(vme_io_vme_wr_0_cmd_valid),
    .io_vme_wr_0_cmd_bits_addr(vme_io_vme_wr_0_cmd_bits_addr),
    .io_vme_wr_0_cmd_bits_len(vme_io_vme_wr_0_cmd_bits_len),
    .io_vme_wr_0_data_ready(vme_io_vme_wr_0_data_ready),
    .io_vme_wr_0_data_valid(vme_io_vme_wr_0_data_valid),
    .io_vme_wr_0_data_bits(vme_io_vme_wr_0_data_bits),
    .io_vme_wr_0_ack(vme_io_vme_wr_0_ack)
  );
  Core core ( // @[VTAShell.scala 50:20:@25003.4]
    .clock(core_clock),
    .reset(core_reset),
    .io_vcr_launch(core_io_vcr_launch),
    .io_vcr_finish(core_io_vcr_finish),
    .io_vcr_ecnt_0_valid(core_io_vcr_ecnt_0_valid),
    .io_vcr_ecnt_0_bits(core_io_vcr_ecnt_0_bits),
    .io_vcr_vals_0(core_io_vcr_vals_0),
    .io_vcr_ptrs_0(core_io_vcr_ptrs_0),
    .io_vcr_ptrs_1(core_io_vcr_ptrs_1),
    .io_vcr_ptrs_2(core_io_vcr_ptrs_2),
    .io_vcr_ptrs_3(core_io_vcr_ptrs_3),
    .io_vcr_ptrs_4(core_io_vcr_ptrs_4),
    .io_vcr_ptrs_5(core_io_vcr_ptrs_5),
    .io_vcr_ucnt_0_valid(core_io_vcr_ucnt_0_valid),
    .io_vcr_ucnt_0_bits(core_io_vcr_ucnt_0_bits),
    .io_vme_rd_0_cmd_ready(core_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(core_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(core_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(core_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(core_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(core_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits(core_io_vme_rd_0_data_bits),
    .io_vme_rd_1_cmd_ready(core_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(core_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(core_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(core_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_data_ready(core_io_vme_rd_1_data_ready),
    .io_vme_rd_1_data_valid(core_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits(core_io_vme_rd_1_data_bits),
    .io_vme_rd_2_cmd_ready(core_io_vme_rd_2_cmd_ready),
    .io_vme_rd_2_cmd_valid(core_io_vme_rd_2_cmd_valid),
    .io_vme_rd_2_cmd_bits_addr(core_io_vme_rd_2_cmd_bits_addr),
    .io_vme_rd_2_cmd_bits_len(core_io_vme_rd_2_cmd_bits_len),
    .io_vme_rd_2_data_ready(core_io_vme_rd_2_data_ready),
    .io_vme_rd_2_data_valid(core_io_vme_rd_2_data_valid),
    .io_vme_rd_2_data_bits(core_io_vme_rd_2_data_bits),
    .io_vme_rd_3_cmd_ready(core_io_vme_rd_3_cmd_ready),
    .io_vme_rd_3_cmd_valid(core_io_vme_rd_3_cmd_valid),
    .io_vme_rd_3_cmd_bits_addr(core_io_vme_rd_3_cmd_bits_addr),
    .io_vme_rd_3_cmd_bits_len(core_io_vme_rd_3_cmd_bits_len),
    .io_vme_rd_3_data_ready(core_io_vme_rd_3_data_ready),
    .io_vme_rd_3_data_valid(core_io_vme_rd_3_data_valid),
    .io_vme_rd_3_data_bits(core_io_vme_rd_3_data_bits),
    .io_vme_rd_4_cmd_ready(core_io_vme_rd_4_cmd_ready),
    .io_vme_rd_4_cmd_valid(core_io_vme_rd_4_cmd_valid),
    .io_vme_rd_4_cmd_bits_addr(core_io_vme_rd_4_cmd_bits_addr),
    .io_vme_rd_4_cmd_bits_len(core_io_vme_rd_4_cmd_bits_len),
    .io_vme_rd_4_data_ready(core_io_vme_rd_4_data_ready),
    .io_vme_rd_4_data_valid(core_io_vme_rd_4_data_valid),
    .io_vme_rd_4_data_bits(core_io_vme_rd_4_data_bits),
    .io_vme_wr_0_cmd_ready(core_io_vme_wr_0_cmd_ready),
    .io_vme_wr_0_cmd_valid(core_io_vme_wr_0_cmd_valid),
    .io_vme_wr_0_cmd_bits_addr(core_io_vme_wr_0_cmd_bits_addr),
    .io_vme_wr_0_cmd_bits_len(core_io_vme_wr_0_cmd_bits_len),
    .io_vme_wr_0_data_ready(core_io_vme_wr_0_data_ready),
    .io_vme_wr_0_data_valid(core_io_vme_wr_0_data_valid),
    .io_vme_wr_0_data_bits(core_io_vme_wr_0_data_bits),
    .io_vme_wr_0_ack(core_io_vme_wr_0_ack)
  );
  assign io_host_aw_ready = vcr_io_host_aw_ready; // @[VTAShell.scala 55:15:@25078.4]
  assign io_host_w_ready = vcr_io_host_w_ready; // @[VTAShell.scala 55:15:@25075.4]
  assign io_host_b_valid = vcr_io_host_b_valid; // @[VTAShell.scala 55:15:@25070.4]
  assign io_host_ar_ready = vcr_io_host_ar_ready; // @[VTAShell.scala 55:15:@25068.4]
  assign io_host_r_valid = vcr_io_host_r_valid; // @[VTAShell.scala 55:15:@25064.4]
  assign io_host_r_bits_data = vcr_io_host_r_bits_data; // @[VTAShell.scala 55:15:@25063.4]
  assign io_mem_aw_valid = vme_io_mem_aw_valid; // @[VTAShell.scala 56:10:@25122.4]
  assign io_mem_aw_bits_addr = vme_io_mem_aw_bits_addr; // @[VTAShell.scala 56:10:@25121.4]
  assign io_mem_aw_bits_len = vme_io_mem_aw_bits_len; // @[VTAShell.scala 56:10:@25118.4]
  assign io_mem_w_valid = vme_io_mem_w_valid; // @[VTAShell.scala 56:10:@25109.4]
  assign io_mem_w_bits_data = vme_io_mem_w_bits_data; // @[VTAShell.scala 56:10:@25108.4]
  assign io_mem_w_bits_last = vme_io_mem_w_bits_last; // @[VTAShell.scala 56:10:@25106.4]
  assign io_mem_ar_valid = vme_io_mem_ar_valid; // @[VTAShell.scala 56:10:@25097.4]
  assign io_mem_ar_bits_addr = vme_io_mem_ar_bits_addr; // @[VTAShell.scala 56:10:@25096.4]
  assign io_mem_ar_bits_len = vme_io_mem_ar_bits_len; // @[VTAShell.scala 56:10:@25093.4]
  assign io_mem_r_ready = vme_io_mem_r_ready; // @[VTAShell.scala 56:10:@25085.4]
  assign vcr_clock = clock; // @[:@24998.4]
  assign vcr_reset = reset; // @[:@24999.4]
  assign vcr_io_host_aw_valid = io_host_aw_valid; // @[VTAShell.scala 55:15:@25077.4]
  assign vcr_io_host_aw_bits_addr = io_host_aw_bits_addr; // @[VTAShell.scala 55:15:@25076.4]
  assign vcr_io_host_w_valid = io_host_w_valid; // @[VTAShell.scala 55:15:@25074.4]
  assign vcr_io_host_w_bits_data = io_host_w_bits_data; // @[VTAShell.scala 55:15:@25073.4]
  assign vcr_io_host_b_ready = io_host_b_ready; // @[VTAShell.scala 55:15:@25071.4]
  assign vcr_io_host_ar_valid = io_host_ar_valid; // @[VTAShell.scala 55:15:@25067.4]
  assign vcr_io_host_ar_bits_addr = io_host_ar_bits_addr; // @[VTAShell.scala 55:15:@25066.4]
  assign vcr_io_host_r_ready = io_host_r_ready; // @[VTAShell.scala 55:15:@25065.4]
  assign vcr_io_vcr_finish = core_io_vcr_finish; // @[VTAShell.scala 52:15:@25017.4]
  assign vcr_io_vcr_ecnt_0_valid = core_io_vcr_ecnt_0_valid; // @[VTAShell.scala 52:15:@25016.4]
  assign vcr_io_vcr_ecnt_0_bits = core_io_vcr_ecnt_0_bits; // @[VTAShell.scala 52:15:@25015.4]
  assign vcr_io_vcr_ucnt_0_valid = core_io_vcr_ucnt_0_valid; // @[VTAShell.scala 52:15:@25007.4]
  assign vcr_io_vcr_ucnt_0_bits = core_io_vcr_ucnt_0_bits; // @[VTAShell.scala 52:15:@25006.4]
  assign vme_clock = clock; // @[:@25001.4]
  assign vme_reset = reset; // @[:@25002.4]
  assign vme_io_mem_aw_ready = io_mem_aw_ready; // @[VTAShell.scala 56:10:@25123.4]
  assign vme_io_mem_w_ready = io_mem_w_ready; // @[VTAShell.scala 56:10:@25110.4]
  assign vme_io_mem_b_valid = io_mem_b_valid; // @[VTAShell.scala 56:10:@25102.4]
  assign vme_io_mem_ar_ready = io_mem_ar_ready; // @[VTAShell.scala 56:10:@25098.4]
  assign vme_io_mem_r_valid = io_mem_r_valid; // @[VTAShell.scala 56:10:@25084.4]
  assign vme_io_mem_r_bits_data = io_mem_r_bits_data; // @[VTAShell.scala 56:10:@25083.4]
  assign vme_io_mem_r_bits_last = io_mem_r_bits_last; // @[VTAShell.scala 56:10:@25081.4]
  assign vme_io_vme_rd_0_cmd_valid = core_io_vme_rd_0_cmd_valid; // @[VTAShell.scala 53:14:@25032.4]
  assign vme_io_vme_rd_0_cmd_bits_addr = core_io_vme_rd_0_cmd_bits_addr; // @[VTAShell.scala 53:14:@25031.4]
  assign vme_io_vme_rd_0_cmd_bits_len = core_io_vme_rd_0_cmd_bits_len; // @[VTAShell.scala 53:14:@25030.4]
  assign vme_io_vme_rd_0_data_ready = core_io_vme_rd_0_data_ready; // @[VTAShell.scala 53:14:@25029.4]
  assign vme_io_vme_rd_1_cmd_valid = core_io_vme_rd_1_cmd_valid; // @[VTAShell.scala 53:14:@25039.4]
  assign vme_io_vme_rd_1_cmd_bits_addr = core_io_vme_rd_1_cmd_bits_addr; // @[VTAShell.scala 53:14:@25038.4]
  assign vme_io_vme_rd_1_cmd_bits_len = core_io_vme_rd_1_cmd_bits_len; // @[VTAShell.scala 53:14:@25037.4]
  assign vme_io_vme_rd_1_data_ready = core_io_vme_rd_1_data_ready; // @[VTAShell.scala 53:14:@25036.4]
  assign vme_io_vme_rd_2_cmd_valid = core_io_vme_rd_2_cmd_valid; // @[VTAShell.scala 53:14:@25046.4]
  assign vme_io_vme_rd_2_cmd_bits_addr = core_io_vme_rd_2_cmd_bits_addr; // @[VTAShell.scala 53:14:@25045.4]
  assign vme_io_vme_rd_2_cmd_bits_len = core_io_vme_rd_2_cmd_bits_len; // @[VTAShell.scala 53:14:@25044.4]
  assign vme_io_vme_rd_2_data_ready = core_io_vme_rd_2_data_ready; // @[VTAShell.scala 53:14:@25043.4]
  assign vme_io_vme_rd_3_cmd_valid = core_io_vme_rd_3_cmd_valid; // @[VTAShell.scala 53:14:@25053.4]
  assign vme_io_vme_rd_3_cmd_bits_addr = core_io_vme_rd_3_cmd_bits_addr; // @[VTAShell.scala 53:14:@25052.4]
  assign vme_io_vme_rd_3_cmd_bits_len = core_io_vme_rd_3_cmd_bits_len; // @[VTAShell.scala 53:14:@25051.4]
  assign vme_io_vme_rd_3_data_ready = core_io_vme_rd_3_data_ready; // @[VTAShell.scala 53:14:@25050.4]
  assign vme_io_vme_rd_4_cmd_valid = core_io_vme_rd_4_cmd_valid; // @[VTAShell.scala 53:14:@25060.4]
  assign vme_io_vme_rd_4_cmd_bits_addr = core_io_vme_rd_4_cmd_bits_addr; // @[VTAShell.scala 53:14:@25059.4]
  assign vme_io_vme_rd_4_cmd_bits_len = core_io_vme_rd_4_cmd_bits_len; // @[VTAShell.scala 53:14:@25058.4]
  assign vme_io_vme_rd_4_data_ready = core_io_vme_rd_4_data_ready; // @[VTAShell.scala 53:14:@25057.4]
  assign vme_io_vme_wr_0_cmd_valid = core_io_vme_wr_0_cmd_valid; // @[VTAShell.scala 53:14:@25025.4]
  assign vme_io_vme_wr_0_cmd_bits_addr = core_io_vme_wr_0_cmd_bits_addr; // @[VTAShell.scala 53:14:@25024.4]
  assign vme_io_vme_wr_0_cmd_bits_len = core_io_vme_wr_0_cmd_bits_len; // @[VTAShell.scala 53:14:@25023.4]
  assign vme_io_vme_wr_0_data_valid = core_io_vme_wr_0_data_valid; // @[VTAShell.scala 53:14:@25021.4]
  assign vme_io_vme_wr_0_data_bits = core_io_vme_wr_0_data_bits; // @[VTAShell.scala 53:14:@25020.4]
  assign core_clock = clock; // @[:@25004.4]
  assign core_reset = reset; // @[:@25005.4]
  assign core_io_vcr_launch = vcr_io_vcr_launch; // @[VTAShell.scala 52:15:@25018.4]
  assign core_io_vcr_vals_0 = vcr_io_vcr_vals_0; // @[VTAShell.scala 52:15:@25014.4]
  assign core_io_vcr_ptrs_0 = vcr_io_vcr_ptrs_0; // @[VTAShell.scala 52:15:@25008.4]
  assign core_io_vcr_ptrs_1 = vcr_io_vcr_ptrs_1; // @[VTAShell.scala 52:15:@25009.4]
  assign core_io_vcr_ptrs_2 = vcr_io_vcr_ptrs_2; // @[VTAShell.scala 52:15:@25010.4]
  assign core_io_vcr_ptrs_3 = vcr_io_vcr_ptrs_3; // @[VTAShell.scala 52:15:@25011.4]
  assign core_io_vcr_ptrs_4 = vcr_io_vcr_ptrs_4; // @[VTAShell.scala 52:15:@25012.4]
  assign core_io_vcr_ptrs_5 = vcr_io_vcr_ptrs_5; // @[VTAShell.scala 52:15:@25013.4]
  assign core_io_vme_rd_0_cmd_ready = vme_io_vme_rd_0_cmd_ready; // @[VTAShell.scala 53:14:@25033.4]
  assign core_io_vme_rd_0_data_valid = vme_io_vme_rd_0_data_valid; // @[VTAShell.scala 53:14:@25028.4]
  assign core_io_vme_rd_0_data_bits = vme_io_vme_rd_0_data_bits; // @[VTAShell.scala 53:14:@25027.4]
  assign core_io_vme_rd_1_cmd_ready = vme_io_vme_rd_1_cmd_ready; // @[VTAShell.scala 53:14:@25040.4]
  assign core_io_vme_rd_1_data_valid = vme_io_vme_rd_1_data_valid; // @[VTAShell.scala 53:14:@25035.4]
  assign core_io_vme_rd_1_data_bits = vme_io_vme_rd_1_data_bits; // @[VTAShell.scala 53:14:@25034.4]
  assign core_io_vme_rd_2_cmd_ready = vme_io_vme_rd_2_cmd_ready; // @[VTAShell.scala 53:14:@25047.4]
  assign core_io_vme_rd_2_data_valid = vme_io_vme_rd_2_data_valid; // @[VTAShell.scala 53:14:@25042.4]
  assign core_io_vme_rd_2_data_bits = vme_io_vme_rd_2_data_bits; // @[VTAShell.scala 53:14:@25041.4]
  assign core_io_vme_rd_3_cmd_ready = vme_io_vme_rd_3_cmd_ready; // @[VTAShell.scala 53:14:@25054.4]
  assign core_io_vme_rd_3_data_valid = vme_io_vme_rd_3_data_valid; // @[VTAShell.scala 53:14:@25049.4]
  assign core_io_vme_rd_3_data_bits = vme_io_vme_rd_3_data_bits; // @[VTAShell.scala 53:14:@25048.4]
  assign core_io_vme_rd_4_cmd_ready = vme_io_vme_rd_4_cmd_ready; // @[VTAShell.scala 53:14:@25061.4]
  assign core_io_vme_rd_4_data_valid = vme_io_vme_rd_4_data_valid; // @[VTAShell.scala 53:14:@25056.4]
  assign core_io_vme_rd_4_data_bits = vme_io_vme_rd_4_data_bits; // @[VTAShell.scala 53:14:@25055.4]
  assign core_io_vme_wr_0_cmd_ready = vme_io_vme_wr_0_cmd_ready; // @[VTAShell.scala 53:14:@25026.4]
  assign core_io_vme_wr_0_data_ready = vme_io_vme_wr_0_data_ready; // @[VTAShell.scala 53:14:@25022.4]
  assign core_io_vme_wr_0_ack = vme_io_vme_wr_0_ack; // @[VTAShell.scala 53:14:@25019.4]
endmodule
module XilinxShell( // @[:@25125.2]
  input         ap_clk, // @[:@25126.4]
  input         ap_rst_n, // @[:@25127.4]
  output        m_axi_gmem_AWVALID, // @[:@25128.4]
  input         m_axi_gmem_AWREADY, // @[:@25128.4]
  output [31:0] m_axi_gmem_AWADDR, // @[:@25128.4]
  output        m_axi_gmem_AWID, // @[:@25128.4]
  output        m_axi_gmem_AWUSER, // @[:@25128.4]
  output [7:0]  m_axi_gmem_AWLEN, // @[:@25128.4]
  output [2:0]  m_axi_gmem_AWSIZE, // @[:@25128.4]
  output [1:0]  m_axi_gmem_AWBURST, // @[:@25128.4]
  output [1:0]  m_axi_gmem_AWLOCK, // @[:@25128.4]
  output [3:0]  m_axi_gmem_AWCACHE, // @[:@25128.4]
  output [2:0]  m_axi_gmem_AWPROT, // @[:@25128.4]
  output [3:0]  m_axi_gmem_AWQOS, // @[:@25128.4]
  output [3:0]  m_axi_gmem_AWREGION, // @[:@25128.4]
  output        m_axi_gmem_WVALID, // @[:@25128.4]
  input         m_axi_gmem_WREADY, // @[:@25128.4]
  output [63:0] m_axi_gmem_WDATA, // @[:@25128.4]
  output [7:0]  m_axi_gmem_WSTRB, // @[:@25128.4]
  output        m_axi_gmem_WLAST, // @[:@25128.4]
  output        m_axi_gmem_WID, // @[:@25128.4]
  output        m_axi_gmem_WUSER, // @[:@25128.4]
  input         m_axi_gmem_BVALID, // @[:@25128.4]
  output        m_axi_gmem_BREADY, // @[:@25128.4]
  input  [1:0]  m_axi_gmem_BRESP, // @[:@25128.4]
  input         m_axi_gmem_BID, // @[:@25128.4]
  input         m_axi_gmem_BUSER, // @[:@25128.4]
  output        m_axi_gmem_ARVALID, // @[:@25128.4]
  input         m_axi_gmem_ARREADY, // @[:@25128.4]
  output [31:0] m_axi_gmem_ARADDR, // @[:@25128.4]
  output        m_axi_gmem_ARID, // @[:@25128.4]
  output        m_axi_gmem_ARUSER, // @[:@25128.4]
  output [7:0]  m_axi_gmem_ARLEN, // @[:@25128.4]
  output [2:0]  m_axi_gmem_ARSIZE, // @[:@25128.4]
  output [1:0]  m_axi_gmem_ARBURST, // @[:@25128.4]
  output [1:0]  m_axi_gmem_ARLOCK, // @[:@25128.4]
  output [3:0]  m_axi_gmem_ARCACHE, // @[:@25128.4]
  output [2:0]  m_axi_gmem_ARPROT, // @[:@25128.4]
  output [3:0]  m_axi_gmem_ARQOS, // @[:@25128.4]
  output [3:0]  m_axi_gmem_ARREGION, // @[:@25128.4]
  input         m_axi_gmem_RVALID, // @[:@25128.4]
  output        m_axi_gmem_RREADY, // @[:@25128.4]
  input  [63:0] m_axi_gmem_RDATA, // @[:@25128.4]
  input  [1:0]  m_axi_gmem_RRESP, // @[:@25128.4]
  input         m_axi_gmem_RLAST, // @[:@25128.4]
  input         m_axi_gmem_RID, // @[:@25128.4]
  input         m_axi_gmem_RUSER, // @[:@25128.4]
  input         s_axi_control_AWVALID, // @[:@25129.4]
  output        s_axi_control_AWREADY, // @[:@25129.4]
  input  [15:0] s_axi_control_AWADDR, // @[:@25129.4]
  input         s_axi_control_WVALID, // @[:@25129.4]
  output        s_axi_control_WREADY, // @[:@25129.4]
  input  [31:0] s_axi_control_WDATA, // @[:@25129.4]
  input  [3:0]  s_axi_control_WSTRB, // @[:@25129.4]
  output        s_axi_control_BVALID, // @[:@25129.4]
  input         s_axi_control_BREADY, // @[:@25129.4]
  output [1:0]  s_axi_control_BRESP, // @[:@25129.4]
  input         s_axi_control_ARVALID, // @[:@25129.4]
  output        s_axi_control_ARREADY, // @[:@25129.4]
  input  [15:0] s_axi_control_ARADDR, // @[:@25129.4]
  output        s_axi_control_RVALID, // @[:@25129.4]
  input         s_axi_control_RREADY, // @[:@25129.4]
  output [31:0] s_axi_control_RDATA, // @[:@25129.4]
  output [1:0]  s_axi_control_RRESP // @[:@25129.4]
);
  wire  shell_clock; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_reset; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_aw_ready; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_aw_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire [15:0] shell_io_host_aw_bits_addr; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_w_ready; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_w_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire [31:0] shell_io_host_w_bits_data; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_b_ready; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_b_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_ar_ready; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_ar_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire [15:0] shell_io_host_ar_bits_addr; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_r_ready; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_host_r_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire [31:0] shell_io_host_r_bits_data; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_aw_ready; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_aw_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire [31:0] shell_io_mem_aw_bits_addr; // @[XilinxShell.scala 43:11:@25132.4]
  wire [7:0] shell_io_mem_aw_bits_len; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_w_ready; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_w_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire [63:0] shell_io_mem_w_bits_data; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_w_bits_last; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_b_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_ar_ready; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_ar_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire [31:0] shell_io_mem_ar_bits_addr; // @[XilinxShell.scala 43:11:@25132.4]
  wire [7:0] shell_io_mem_ar_bits_len; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_r_ready; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_r_valid; // @[XilinxShell.scala 43:11:@25132.4]
  wire [63:0] shell_io_mem_r_bits_data; // @[XilinxShell.scala 43:11:@25132.4]
  wire  shell_io_mem_r_bits_last; // @[XilinxShell.scala 43:11:@25132.4]
  VTAShell shell ( // @[XilinxShell.scala 43:11:@25132.4]
    .clock(shell_clock),
    .reset(shell_reset),
    .io_host_aw_ready(shell_io_host_aw_ready),
    .io_host_aw_valid(shell_io_host_aw_valid),
    .io_host_aw_bits_addr(shell_io_host_aw_bits_addr),
    .io_host_w_ready(shell_io_host_w_ready),
    .io_host_w_valid(shell_io_host_w_valid),
    .io_host_w_bits_data(shell_io_host_w_bits_data),
    .io_host_b_ready(shell_io_host_b_ready),
    .io_host_b_valid(shell_io_host_b_valid),
    .io_host_ar_ready(shell_io_host_ar_ready),
    .io_host_ar_valid(shell_io_host_ar_valid),
    .io_host_ar_bits_addr(shell_io_host_ar_bits_addr),
    .io_host_r_ready(shell_io_host_r_ready),
    .io_host_r_valid(shell_io_host_r_valid),
    .io_host_r_bits_data(shell_io_host_r_bits_data),
    .io_mem_aw_ready(shell_io_mem_aw_ready),
    .io_mem_aw_valid(shell_io_mem_aw_valid),
    .io_mem_aw_bits_addr(shell_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(shell_io_mem_aw_bits_len),
    .io_mem_w_ready(shell_io_mem_w_ready),
    .io_mem_w_valid(shell_io_mem_w_valid),
    .io_mem_w_bits_data(shell_io_mem_w_bits_data),
    .io_mem_w_bits_last(shell_io_mem_w_bits_last),
    .io_mem_b_valid(shell_io_mem_b_valid),
    .io_mem_ar_ready(shell_io_mem_ar_ready),
    .io_mem_ar_valid(shell_io_mem_ar_valid),
    .io_mem_ar_bits_addr(shell_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(shell_io_mem_ar_bits_len),
    .io_mem_r_ready(shell_io_mem_r_ready),
    .io_mem_r_valid(shell_io_mem_r_valid),
    .io_mem_r_bits_data(shell_io_mem_r_bits_data),
    .io_mem_r_bits_last(shell_io_mem_r_bits_last)
  );
  assign m_axi_gmem_AWVALID = shell_io_mem_aw_valid; // @[XilinxShell.scala 47:22:@25135.4]
  assign m_axi_gmem_AWADDR = shell_io_mem_aw_bits_addr; // @[XilinxShell.scala 49:21:@25137.4]
  assign m_axi_gmem_AWID = 1'h0; // @[XilinxShell.scala 50:19:@25138.4]
  assign m_axi_gmem_AWUSER = 1'h1; // @[XilinxShell.scala 51:21:@25139.4]
  assign m_axi_gmem_AWLEN = shell_io_mem_aw_bits_len; // @[XilinxShell.scala 52:20:@25140.4]
  assign m_axi_gmem_AWSIZE = 3'h3; // @[XilinxShell.scala 53:21:@25141.4]
  assign m_axi_gmem_AWBURST = 2'h1; // @[XilinxShell.scala 54:22:@25142.4]
  assign m_axi_gmem_AWLOCK = 2'h0; // @[XilinxShell.scala 55:21:@25143.4]
  assign m_axi_gmem_AWCACHE = 4'hf; // @[XilinxShell.scala 56:22:@25144.4]
  assign m_axi_gmem_AWPROT = 3'h4; // @[XilinxShell.scala 57:21:@25145.4]
  assign m_axi_gmem_AWQOS = 4'h0; // @[XilinxShell.scala 58:20:@25146.4]
  assign m_axi_gmem_AWREGION = 4'h0; // @[XilinxShell.scala 59:23:@25147.4]
  assign m_axi_gmem_WVALID = shell_io_mem_w_valid; // @[XilinxShell.scala 61:21:@25148.4]
  assign m_axi_gmem_WDATA = shell_io_mem_w_bits_data; // @[XilinxShell.scala 63:20:@25150.4]
  assign m_axi_gmem_WSTRB = 8'hff; // @[XilinxShell.scala 64:20:@25151.4]
  assign m_axi_gmem_WLAST = shell_io_mem_w_bits_last; // @[XilinxShell.scala 65:20:@25152.4]
  assign m_axi_gmem_WID = 1'h0; // @[XilinxShell.scala 66:18:@25153.4]
  assign m_axi_gmem_WUSER = 1'h1; // @[XilinxShell.scala 67:20:@25154.4]
  assign m_axi_gmem_BREADY = shell_io_mem_b_valid; // @[XilinxShell.scala 70:21:@25156.4]
  assign m_axi_gmem_ARVALID = shell_io_mem_ar_valid; // @[XilinxShell.scala 75:22:@25160.4]
  assign m_axi_gmem_ARADDR = shell_io_mem_ar_bits_addr; // @[XilinxShell.scala 77:21:@25162.4]
  assign m_axi_gmem_ARID = 1'h0; // @[XilinxShell.scala 78:19:@25163.4]
  assign m_axi_gmem_ARUSER = 1'h1; // @[XilinxShell.scala 79:21:@25164.4]
  assign m_axi_gmem_ARLEN = shell_io_mem_ar_bits_len; // @[XilinxShell.scala 80:20:@25165.4]
  assign m_axi_gmem_ARSIZE = 3'h3; // @[XilinxShell.scala 81:21:@25166.4]
  assign m_axi_gmem_ARBURST = 2'h1; // @[XilinxShell.scala 82:22:@25167.4]
  assign m_axi_gmem_ARLOCK = 2'h0; // @[XilinxShell.scala 83:21:@25168.4]
  assign m_axi_gmem_ARCACHE = 4'hf; // @[XilinxShell.scala 84:22:@25169.4]
  assign m_axi_gmem_ARPROT = 3'h4; // @[XilinxShell.scala 85:21:@25170.4]
  assign m_axi_gmem_ARQOS = 4'h0; // @[XilinxShell.scala 86:20:@25171.4]
  assign m_axi_gmem_ARREGION = 4'h0; // @[XilinxShell.scala 87:23:@25172.4]
  assign m_axi_gmem_RREADY = shell_io_mem_r_ready; // @[XilinxShell.scala 90:21:@25174.4]
  assign s_axi_control_AWREADY = shell_io_host_aw_ready; // @[XilinxShell.scala 99:25:@25181.4]
  assign s_axi_control_WREADY = shell_io_host_w_ready; // @[XilinxShell.scala 103:24:@25184.4]
  assign s_axi_control_BVALID = shell_io_host_b_valid; // @[XilinxShell.scala 107:24:@25187.4]
  assign s_axi_control_BRESP = 2'h0; // @[XilinxShell.scala 109:23:@25189.4]
  assign s_axi_control_ARREADY = shell_io_host_ar_ready; // @[XilinxShell.scala 112:25:@25191.4]
  assign s_axi_control_RVALID = shell_io_host_r_valid; // @[XilinxShell.scala 115:24:@25193.4]
  assign s_axi_control_RDATA = shell_io_host_r_bits_data; // @[XilinxShell.scala 117:23:@25195.4]
  assign s_axi_control_RRESP = 2'h0; // @[XilinxShell.scala 118:23:@25196.4]
  assign shell_clock = ap_clk; // @[:@25133.4]
  assign shell_reset = ~ ap_rst_n; // @[:@25134.4]
  assign shell_io_host_aw_valid = s_axi_control_AWVALID; // @[XilinxShell.scala 98:26:@25180.4]
  assign shell_io_host_aw_bits_addr = s_axi_control_AWADDR; // @[XilinxShell.scala 100:30:@25182.4]
  assign shell_io_host_w_valid = s_axi_control_WVALID; // @[XilinxShell.scala 102:25:@25183.4]
  assign shell_io_host_w_bits_data = s_axi_control_WDATA; // @[XilinxShell.scala 104:29:@25185.4]
  assign shell_io_host_b_ready = s_axi_control_BREADY; // @[XilinxShell.scala 108:25:@25188.4]
  assign shell_io_host_ar_valid = s_axi_control_ARVALID; // @[XilinxShell.scala 111:26:@25190.4]
  assign shell_io_host_ar_bits_addr = s_axi_control_ARADDR; // @[XilinxShell.scala 113:30:@25192.4]
  assign shell_io_host_r_ready = s_axi_control_RREADY; // @[XilinxShell.scala 116:25:@25194.4]
  assign shell_io_mem_aw_ready = m_axi_gmem_AWREADY; // @[XilinxShell.scala 48:25:@25136.4]
  assign shell_io_mem_w_ready = m_axi_gmem_WREADY; // @[XilinxShell.scala 62:24:@25149.4]
  assign shell_io_mem_b_valid = m_axi_gmem_BVALID; // @[XilinxShell.scala 69:24:@25155.4]
  assign shell_io_mem_ar_ready = m_axi_gmem_ARREADY; // @[XilinxShell.scala 76:25:@25161.4]
  assign shell_io_mem_r_valid = m_axi_gmem_RVALID; // @[XilinxShell.scala 89:24:@25173.4]
  assign shell_io_mem_r_bits_data = m_axi_gmem_RDATA; // @[XilinxShell.scala 91:28:@25175.4]
  assign shell_io_mem_r_bits_last = m_axi_gmem_RLAST; // @[XilinxShell.scala 93:28:@25177.4]
endmodule
