module VTASim( // @[:@11.2]
  input   clock, // @[:@12.4]
  input   reset, // @[:@13.4]
  output  sim_wait // @[:@14.4]
);
  wire  sim_dpi_wait; // @[SimShell.scala 74:19:@16.4]
  wire  sim_reset; // @[SimShell.scala 74:19:@16.4]
  wire  sim_clock; // @[SimShell.scala 74:19:@16.4]
  VTASimDPI sim ( // @[SimShell.scala 74:19:@16.4]
    .dpi_wait(sim_dpi_wait),
    .reset(sim_reset),
    .clock(sim_clock)
  );
  assign sim_wait = sim_dpi_wait; // @[SimShell.scala 77:12:@22.4]
  assign sim_reset = reset; // @[SimShell.scala 75:16:@20.4]
  assign sim_clock = clock; // @[SimShell.scala 76:16:@21.4]
endmodule
module VTAHostDPIToAXI( // @[:@32.2]
  input         clock, // @[:@33.4]
  input         reset, // @[:@34.4]
  input         io_dpi_req_valid, // @[:@35.4]
  input         io_dpi_req_opcode, // @[:@35.4]
  input  [7:0]  io_dpi_req_addr, // @[:@35.4]
  input  [31:0] io_dpi_req_value, // @[:@35.4]
  output        io_dpi_req_deq, // @[:@35.4]
  output        io_dpi_resp_valid, // @[:@35.4]
  output [31:0] io_dpi_resp_bits, // @[:@35.4]
  input         io_axi_aw_ready, // @[:@35.4]
  output        io_axi_aw_valid, // @[:@35.4]
  output [15:0] io_axi_aw_bits_addr, // @[:@35.4]
  input         io_axi_w_ready, // @[:@35.4]
  output        io_axi_w_valid, // @[:@35.4]
  output [31:0] io_axi_w_bits_data, // @[:@35.4]
  output        io_axi_b_ready, // @[:@35.4]
  input         io_axi_b_valid, // @[:@35.4]
  input         io_axi_ar_ready, // @[:@35.4]
  output        io_axi_ar_valid, // @[:@35.4]
  output [15:0] io_axi_ar_bits_addr, // @[:@35.4]
  output        io_axi_r_ready, // @[:@35.4]
  input         io_axi_r_valid, // @[:@35.4]
  input  [31:0] io_axi_r_bits_data // @[:@35.4]
);
  reg [7:0] addr; // @[VTAHostDPI.scala 86:21:@39.4]
  reg [31:0] _RAND_0;
  reg [31:0] data; // @[VTAHostDPI.scala 87:21:@42.4]
  reg [31:0] _RAND_1;
  reg [2:0] state; // @[VTAHostDPI.scala 90:22:@43.4]
  reg [31:0] _RAND_2;
  wire  _T_72; // @[Conditional.scala 37:30:@44.4]
  wire [2:0] _GEN_0; // @[VTAHostDPI.scala 95:33:@47.8]
  wire [2:0] _GEN_1; // @[VTAHostDPI.scala 94:30:@46.6]
  wire  _T_73; // @[Conditional.scala 37:30:@56.6]
  wire [2:0] _GEN_2; // @[VTAHostDPI.scala 103:29:@58.8]
  wire  _T_74; // @[Conditional.scala 37:30:@63.8]
  wire [2:0] _GEN_3; // @[VTAHostDPI.scala 108:28:@65.10]
  wire  _T_75; // @[Conditional.scala 37:30:@70.10]
  wire [2:0] _GEN_4; // @[VTAHostDPI.scala 113:29:@72.12]
  wire  _T_76; // @[Conditional.scala 37:30:@77.12]
  wire [2:0] _GEN_5; // @[VTAHostDPI.scala 118:28:@79.14]
  wire  _T_77; // @[Conditional.scala 37:30:@84.14]
  wire [2:0] _GEN_6; // @[VTAHostDPI.scala 123:28:@86.16]
  wire [2:0] _GEN_7; // @[Conditional.scala 39:67:@85.14]
  wire [2:0] _GEN_8; // @[Conditional.scala 39:67:@78.12]
  wire [2:0] _GEN_9; // @[Conditional.scala 39:67:@71.10]
  wire [2:0] _GEN_10; // @[Conditional.scala 39:67:@64.8]
  wire [2:0] _GEN_11; // @[Conditional.scala 39:67:@57.6]
  wire [2:0] _GEN_12; // @[Conditional.scala 40:58:@45.4]
  wire  _T_78; // @[VTAHostDPI.scala 129:14:@90.4]
  wire  _T_79; // @[VTAHostDPI.scala 129:24:@91.4]
  wire [7:0] _GEN_13; // @[VTAHostDPI.scala 129:45:@92.4]
  wire [31:0] _GEN_14; // @[VTAHostDPI.scala 129:45:@92.4]
  wire  _T_80; // @[VTAHostDPI.scala 134:28:@96.4]
  wire  _T_84; // @[VTAHostDPI.scala 141:28:@105.4]
  wire  _T_87; // @[VTAHostDPI.scala 145:45:@111.4]
  wire  _T_89; // @[VTAHostDPI.scala 145:91:@113.4]
  assign _T_72 = 3'h0 == state; // @[Conditional.scala 37:30:@44.4]
  assign _GEN_0 = io_dpi_req_opcode ? 3'h3 : 3'h1; // @[VTAHostDPI.scala 95:33:@47.8]
  assign _GEN_1 = io_dpi_req_valid ? _GEN_0 : state; // @[VTAHostDPI.scala 94:30:@46.6]
  assign _T_73 = 3'h1 == state; // @[Conditional.scala 37:30:@56.6]
  assign _GEN_2 = io_axi_ar_ready ? 3'h2 : state; // @[VTAHostDPI.scala 103:29:@58.8]
  assign _T_74 = 3'h2 == state; // @[Conditional.scala 37:30:@63.8]
  assign _GEN_3 = io_axi_r_valid ? 3'h0 : state; // @[VTAHostDPI.scala 108:28:@65.10]
  assign _T_75 = 3'h3 == state; // @[Conditional.scala 37:30:@70.10]
  assign _GEN_4 = io_axi_aw_ready ? 3'h4 : state; // @[VTAHostDPI.scala 113:29:@72.12]
  assign _T_76 = 3'h4 == state; // @[Conditional.scala 37:30:@77.12]
  assign _GEN_5 = io_axi_w_ready ? 3'h5 : state; // @[VTAHostDPI.scala 118:28:@79.14]
  assign _T_77 = 3'h5 == state; // @[Conditional.scala 37:30:@84.14]
  assign _GEN_6 = io_axi_b_valid ? 3'h0 : state; // @[VTAHostDPI.scala 123:28:@86.16]
  assign _GEN_7 = _T_77 ? _GEN_6 : state; // @[Conditional.scala 39:67:@85.14]
  assign _GEN_8 = _T_76 ? _GEN_5 : _GEN_7; // @[Conditional.scala 39:67:@78.12]
  assign _GEN_9 = _T_75 ? _GEN_4 : _GEN_8; // @[Conditional.scala 39:67:@71.10]
  assign _GEN_10 = _T_74 ? _GEN_3 : _GEN_9; // @[Conditional.scala 39:67:@64.8]
  assign _GEN_11 = _T_73 ? _GEN_2 : _GEN_10; // @[Conditional.scala 39:67:@57.6]
  assign _GEN_12 = _T_72 ? _GEN_1 : _GEN_11; // @[Conditional.scala 40:58:@45.4]
  assign _T_78 = state == 3'h0; // @[VTAHostDPI.scala 129:14:@90.4]
  assign _T_79 = _T_78 & io_dpi_req_valid; // @[VTAHostDPI.scala 129:24:@91.4]
  assign _GEN_13 = _T_79 ? io_dpi_req_addr : addr; // @[VTAHostDPI.scala 129:45:@92.4]
  assign _GEN_14 = _T_79 ? io_dpi_req_value : data; // @[VTAHostDPI.scala 129:45:@92.4]
  assign _T_80 = state == 3'h3; // @[VTAHostDPI.scala 134:28:@96.4]
  assign _T_84 = state == 3'h1; // @[VTAHostDPI.scala 141:28:@105.4]
  assign _T_87 = _T_84 & io_axi_ar_ready; // @[VTAHostDPI.scala 145:45:@111.4]
  assign _T_89 = _T_80 & io_axi_aw_ready; // @[VTAHostDPI.scala 145:91:@113.4]
  assign io_dpi_req_deq = _T_87 | _T_89; // @[VTAHostDPI.scala 145:18:@115.4]
  assign io_dpi_resp_valid = io_axi_r_valid; // @[VTAHostDPI.scala 146:21:@116.4]
  assign io_dpi_resp_bits = io_axi_r_bits_data; // @[VTAHostDPI.scala 147:20:@117.4]
  assign io_axi_aw_valid = state == 3'h3; // @[VTAHostDPI.scala 134:19:@97.4]
  assign io_axi_aw_bits_addr = {{8'd0}, addr}; // @[VTAHostDPI.scala 135:23:@98.4]
  assign io_axi_w_valid = state == 3'h4; // @[VTAHostDPI.scala 136:18:@100.4]
  assign io_axi_w_bits_data = data; // @[VTAHostDPI.scala 137:22:@101.4]
  assign io_axi_b_ready = state == 3'h5; // @[VTAHostDPI.scala 139:18:@104.4]
  assign io_axi_ar_valid = state == 3'h1; // @[VTAHostDPI.scala 141:19:@106.4]
  assign io_axi_ar_bits_addr = {{8'd0}, addr}; // @[VTAHostDPI.scala 142:23:@107.4]
  assign io_axi_r_ready = state == 3'h2; // @[VTAHostDPI.scala 143:18:@109.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      addr <= 8'h0;
    end else begin
      if (_T_79) begin
        addr <= io_dpi_req_addr;
      end
    end
    if (reset) begin
      data <= 32'h0;
    end else begin
      if (_T_79) begin
        data <= io_dpi_req_value;
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_72) begin
        if (io_dpi_req_valid) begin
          if (io_dpi_req_opcode) begin
            state <= 3'h3;
          end else begin
            state <= 3'h1;
          end
        end
      end else begin
        if (_T_73) begin
          if (io_axi_ar_ready) begin
            state <= 3'h2;
          end
        end else begin
          if (_T_74) begin
            if (io_axi_r_valid) begin
              state <= 3'h0;
            end
          end else begin
            if (_T_75) begin
              if (io_axi_aw_ready) begin
                state <= 3'h4;
              end
            end else begin
              if (_T_76) begin
                if (io_axi_w_ready) begin
                  state <= 3'h5;
                end
              end else begin
                if (_T_77) begin
                  if (io_axi_b_valid) begin
                    state <= 3'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module VTAHost( // @[:@119.2]
  input         clock, // @[:@120.4]
  input         reset, // @[:@121.4]
  input         io_axi_aw_ready, // @[:@122.4]
  output        io_axi_aw_valid, // @[:@122.4]
  output [15:0] io_axi_aw_bits_addr, // @[:@122.4]
  input         io_axi_w_ready, // @[:@122.4]
  output        io_axi_w_valid, // @[:@122.4]
  output [31:0] io_axi_w_bits_data, // @[:@122.4]
  output        io_axi_b_ready, // @[:@122.4]
  input         io_axi_b_valid, // @[:@122.4]
  input         io_axi_ar_ready, // @[:@122.4]
  output        io_axi_ar_valid, // @[:@122.4]
  output [15:0] io_axi_ar_bits_addr, // @[:@122.4]
  output        io_axi_r_ready, // @[:@122.4]
  input         io_axi_r_valid, // @[:@122.4]
  input  [31:0] io_axi_r_bits_data // @[:@122.4]
);
  wire  host_dpi_dpi_req_valid; // @[SimShell.scala 39:24:@124.4]
  wire  host_dpi_dpi_req_opcode; // @[SimShell.scala 39:24:@124.4]
  wire [7:0] host_dpi_dpi_req_addr; // @[SimShell.scala 39:24:@124.4]
  wire [31:0] host_dpi_dpi_req_value; // @[SimShell.scala 39:24:@124.4]
  wire  host_dpi_dpi_req_deq; // @[SimShell.scala 39:24:@124.4]
  wire  host_dpi_dpi_resp_valid; // @[SimShell.scala 39:24:@124.4]
  wire [31:0] host_dpi_dpi_resp_bits; // @[SimShell.scala 39:24:@124.4]
  wire  host_dpi_reset; // @[SimShell.scala 39:24:@124.4]
  wire  host_dpi_clock; // @[SimShell.scala 39:24:@124.4]
  wire  host_axi_clock; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_reset; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_dpi_req_valid; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_dpi_req_opcode; // @[SimShell.scala 40:24:@128.4]
  wire [7:0] host_axi_io_dpi_req_addr; // @[SimShell.scala 40:24:@128.4]
  wire [31:0] host_axi_io_dpi_req_value; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_dpi_req_deq; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_dpi_resp_valid; // @[SimShell.scala 40:24:@128.4]
  wire [31:0] host_axi_io_dpi_resp_bits; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_aw_ready; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_aw_valid; // @[SimShell.scala 40:24:@128.4]
  wire [15:0] host_axi_io_axi_aw_bits_addr; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_w_ready; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_w_valid; // @[SimShell.scala 40:24:@128.4]
  wire [31:0] host_axi_io_axi_w_bits_data; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_b_ready; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_b_valid; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_ar_ready; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_ar_valid; // @[SimShell.scala 40:24:@128.4]
  wire [15:0] host_axi_io_axi_ar_bits_addr; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_r_ready; // @[SimShell.scala 40:24:@128.4]
  wire  host_axi_io_axi_r_valid; // @[SimShell.scala 40:24:@128.4]
  wire [31:0] host_axi_io_axi_r_bits_data; // @[SimShell.scala 40:24:@128.4]
  VTAHostDPI host_dpi ( // @[SimShell.scala 39:24:@124.4]
    .dpi_req_valid(host_dpi_dpi_req_valid),
    .dpi_req_opcode(host_dpi_dpi_req_opcode),
    .dpi_req_addr(host_dpi_dpi_req_addr),
    .dpi_req_value(host_dpi_dpi_req_value),
    .dpi_req_deq(host_dpi_dpi_req_deq),
    .dpi_resp_valid(host_dpi_dpi_resp_valid),
    .dpi_resp_bits(host_dpi_dpi_resp_bits),
    .reset(host_dpi_reset),
    .clock(host_dpi_clock)
  );
  VTAHostDPIToAXI host_axi ( // @[SimShell.scala 40:24:@128.4]
    .clock(host_axi_clock),
    .reset(host_axi_reset),
    .io_dpi_req_valid(host_axi_io_dpi_req_valid),
    .io_dpi_req_opcode(host_axi_io_dpi_req_opcode),
    .io_dpi_req_addr(host_axi_io_dpi_req_addr),
    .io_dpi_req_value(host_axi_io_dpi_req_value),
    .io_dpi_req_deq(host_axi_io_dpi_req_deq),
    .io_dpi_resp_valid(host_axi_io_dpi_resp_valid),
    .io_dpi_resp_bits(host_axi_io_dpi_resp_bits),
    .io_axi_aw_ready(host_axi_io_axi_aw_ready),
    .io_axi_aw_valid(host_axi_io_axi_aw_valid),
    .io_axi_aw_bits_addr(host_axi_io_axi_aw_bits_addr),
    .io_axi_w_ready(host_axi_io_axi_w_ready),
    .io_axi_w_valid(host_axi_io_axi_w_valid),
    .io_axi_w_bits_data(host_axi_io_axi_w_bits_data),
    .io_axi_b_ready(host_axi_io_axi_b_ready),
    .io_axi_b_valid(host_axi_io_axi_b_valid),
    .io_axi_ar_ready(host_axi_io_axi_ar_ready),
    .io_axi_ar_valid(host_axi_io_axi_ar_valid),
    .io_axi_ar_bits_addr(host_axi_io_axi_ar_bits_addr),
    .io_axi_r_ready(host_axi_io_axi_r_ready),
    .io_axi_r_valid(host_axi_io_axi_r_valid),
    .io_axi_r_bits_data(host_axi_io_axi_r_bits_data)
  );
  assign io_axi_aw_valid = host_axi_io_axi_aw_valid; // @[SimShell.scala 44:10:@155.4]
  assign io_axi_aw_bits_addr = host_axi_io_axi_aw_bits_addr; // @[SimShell.scala 44:10:@154.4]
  assign io_axi_w_valid = host_axi_io_axi_w_valid; // @[SimShell.scala 44:10:@152.4]
  assign io_axi_w_bits_data = host_axi_io_axi_w_bits_data; // @[SimShell.scala 44:10:@151.4]
  assign io_axi_b_ready = host_axi_io_axi_b_ready; // @[SimShell.scala 44:10:@149.4]
  assign io_axi_ar_valid = host_axi_io_axi_ar_valid; // @[SimShell.scala 44:10:@145.4]
  assign io_axi_ar_bits_addr = host_axi_io_axi_ar_bits_addr; // @[SimShell.scala 44:10:@144.4]
  assign io_axi_r_ready = host_axi_io_axi_r_ready; // @[SimShell.scala 44:10:@143.4]
  assign host_dpi_dpi_req_deq = host_axi_io_dpi_req_deq; // @[SimShell.scala 43:19:@135.4]
  assign host_dpi_dpi_resp_valid = host_axi_io_dpi_resp_valid; // @[SimShell.scala 43:19:@134.4]
  assign host_dpi_dpi_resp_bits = host_axi_io_dpi_resp_bits; // @[SimShell.scala 43:19:@133.4]
  assign host_dpi_reset = reset; // @[SimShell.scala 41:21:@131.4]
  assign host_dpi_clock = clock; // @[SimShell.scala 42:21:@132.4]
  assign host_axi_clock = clock; // @[:@129.4]
  assign host_axi_reset = reset; // @[:@130.4]
  assign host_axi_io_dpi_req_valid = host_dpi_dpi_req_valid; // @[SimShell.scala 43:19:@139.4]
  assign host_axi_io_dpi_req_opcode = host_dpi_dpi_req_opcode; // @[SimShell.scala 43:19:@138.4]
  assign host_axi_io_dpi_req_addr = host_dpi_dpi_req_addr; // @[SimShell.scala 43:19:@137.4]
  assign host_axi_io_dpi_req_value = host_dpi_dpi_req_value; // @[SimShell.scala 43:19:@136.4]
  assign host_axi_io_axi_aw_ready = io_axi_aw_ready; // @[SimShell.scala 44:10:@156.4]
  assign host_axi_io_axi_w_ready = io_axi_w_ready; // @[SimShell.scala 44:10:@153.4]
  assign host_axi_io_axi_b_valid = io_axi_b_valid; // @[SimShell.scala 44:10:@148.4]
  assign host_axi_io_axi_ar_ready = io_axi_ar_ready; // @[SimShell.scala 44:10:@146.4]
  assign host_axi_io_axi_r_valid = io_axi_r_valid; // @[SimShell.scala 44:10:@142.4]
  assign host_axi_io_axi_r_bits_data = io_axi_r_bits_data; // @[SimShell.scala 44:10:@141.4]
endmodule
module VTAMemDPIToAXI( // @[:@166.2]
  input         clock, // @[:@167.4]
  input         reset, // @[:@168.4]
  output        io_dpi_req_valid, // @[:@169.4]
  output        io_dpi_req_opcode, // @[:@169.4]
  output [7:0]  io_dpi_req_len, // @[:@169.4]
  output [63:0] io_dpi_req_addr, // @[:@169.4]
  output        io_dpi_wr_valid, // @[:@169.4]
  output [63:0] io_dpi_wr_bits, // @[:@169.4]
  output        io_dpi_rd_ready, // @[:@169.4]
  input         io_dpi_rd_valid, // @[:@169.4]
  input  [63:0] io_dpi_rd_bits, // @[:@169.4]
  output        io_axi_aw_ready, // @[:@169.4]
  input         io_axi_aw_valid, // @[:@169.4]
  input  [31:0] io_axi_aw_bits_addr, // @[:@169.4]
  input  [7:0]  io_axi_aw_bits_len, // @[:@169.4]
  output        io_axi_w_ready, // @[:@169.4]
  input         io_axi_w_valid, // @[:@169.4]
  input  [63:0] io_axi_w_bits_data, // @[:@169.4]
  input         io_axi_w_bits_last, // @[:@169.4]
  input         io_axi_b_ready, // @[:@169.4]
  output        io_axi_b_valid, // @[:@169.4]
  output        io_axi_ar_ready, // @[:@169.4]
  input         io_axi_ar_valid, // @[:@169.4]
  input  [31:0] io_axi_ar_bits_addr, // @[:@169.4]
  input  [7:0]  io_axi_ar_bits_len, // @[:@169.4]
  input         io_axi_r_ready, // @[:@169.4]
  output        io_axi_r_valid, // @[:@169.4]
  output [63:0] io_axi_r_bits_data, // @[:@169.4]
  output        io_axi_r_bits_last // @[:@169.4]
);
  reg  opcode; // @[VTAMemDPI.scala 83:23:@171.4]
  reg [31:0] _RAND_0;
  reg [7:0] len; // @[VTAMemDPI.scala 84:20:@174.4]
  reg [31:0] _RAND_1;
  reg [63:0] addr; // @[VTAMemDPI.scala 85:21:@177.4]
  reg [63:0] _RAND_2;
  reg [2:0] state; // @[VTAMemDPI.scala 88:22:@178.4]
  reg [31:0] _RAND_3;
  wire  _T_90; // @[Conditional.scala 37:30:@179.4]
  wire [2:0] _GEN_0; // @[VTAMemDPI.scala 94:35:@185.8]
  wire [2:0] _GEN_1; // @[VTAMemDPI.scala 92:29:@181.6]
  wire  _T_91; // @[Conditional.scala 37:30:@190.6]
  wire [2:0] _GEN_2; // @[VTAMemDPI.scala 99:29:@192.8]
  wire  _T_92; // @[Conditional.scala 37:30:@197.8]
  wire  _T_93; // @[VTAMemDPI.scala 104:27:@199.10]
  wire  _T_95; // @[VTAMemDPI.scala 104:53:@200.10]
  wire  _T_96; // @[VTAMemDPI.scala 104:46:@201.10]
  wire [2:0] _GEN_3; // @[VTAMemDPI.scala 104:62:@202.10]
  wire  _T_97; // @[Conditional.scala 37:30:@207.10]
  wire [2:0] _GEN_4; // @[VTAMemDPI.scala 109:29:@209.12]
  wire  _T_98; // @[Conditional.scala 37:30:@214.12]
  wire  _T_99; // @[VTAMemDPI.scala 114:27:@216.14]
  wire [2:0] _GEN_5; // @[VTAMemDPI.scala 114:50:@217.14]
  wire  _T_100; // @[Conditional.scala 37:30:@222.14]
  wire [2:0] _GEN_6; // @[VTAMemDPI.scala 119:28:@224.16]
  wire [2:0] _GEN_7; // @[Conditional.scala 39:67:@223.14]
  wire [2:0] _GEN_8; // @[Conditional.scala 39:67:@215.12]
  wire [2:0] _GEN_9; // @[Conditional.scala 39:67:@208.10]
  wire [2:0] _GEN_10; // @[Conditional.scala 39:67:@198.8]
  wire [2:0] _GEN_11; // @[Conditional.scala 39:67:@191.6]
  wire [2:0] _GEN_12; // @[Conditional.scala 40:58:@180.4]
  wire  _T_101; // @[VTAMemDPI.scala 125:14:@228.4]
  wire  _GEN_13; // @[VTAMemDPI.scala 130:33:@236.8]
  wire [7:0] _GEN_14; // @[VTAMemDPI.scala 130:33:@236.8]
  wire [63:0] _GEN_15; // @[VTAMemDPI.scala 130:33:@236.8]
  wire  _GEN_16; // @[VTAMemDPI.scala 126:27:@230.6]
  wire [7:0] _GEN_17; // @[VTAMemDPI.scala 126:27:@230.6]
  wire [63:0] _GEN_18; // @[VTAMemDPI.scala 126:27:@230.6]
  wire  _T_104; // @[VTAMemDPI.scala 135:20:@243.6]
  wire  _T_107; // @[VTAMemDPI.scala 136:51:@246.8]
  wire  _T_108; // @[VTAMemDPI.scala 136:44:@247.8]
  wire [8:0] _T_110; // @[VTAMemDPI.scala 137:18:@249.10]
  wire [8:0] _T_111; // @[VTAMemDPI.scala 137:18:@250.10]
  wire [7:0] _T_112; // @[VTAMemDPI.scala 137:18:@251.10]
  wire [7:0] _GEN_19; // @[VTAMemDPI.scala 136:60:@248.8]
  wire [7:0] _GEN_20; // @[VTAMemDPI.scala 135:35:@244.6]
  wire  _GEN_21; // @[VTAMemDPI.scala 125:25:@229.4]
  wire [7:0] _GEN_22; // @[VTAMemDPI.scala 125:25:@229.4]
  wire [63:0] _GEN_23; // @[VTAMemDPI.scala 125:25:@229.4]
  wire  _T_113; // @[VTAMemDPI.scala 141:30:@255.4]
  wire  _T_114; // @[VTAMemDPI.scala 141:47:@256.4]
  wire  _T_115; // @[VTAMemDPI.scala 141:75:@257.4]
  wire  _T_116; // @[VTAMemDPI.scala 141:93:@258.4]
  wire  _T_129; // @[VTAMemDPI.scala 157:28:@280.4]
  assign _T_90 = 3'h0 == state; // @[Conditional.scala 37:30:@179.4]
  assign _GEN_0 = io_axi_aw_valid ? 3'h3 : state; // @[VTAMemDPI.scala 94:35:@185.8]
  assign _GEN_1 = io_axi_ar_valid ? 3'h1 : _GEN_0; // @[VTAMemDPI.scala 92:29:@181.6]
  assign _T_91 = 3'h1 == state; // @[Conditional.scala 37:30:@190.6]
  assign _GEN_2 = io_axi_ar_valid ? 3'h2 : state; // @[VTAMemDPI.scala 99:29:@192.8]
  assign _T_92 = 3'h2 == state; // @[Conditional.scala 37:30:@197.8]
  assign _T_93 = io_axi_r_ready & io_dpi_rd_valid; // @[VTAMemDPI.scala 104:27:@199.10]
  assign _T_95 = len == 8'h0; // @[VTAMemDPI.scala 104:53:@200.10]
  assign _T_96 = _T_93 & _T_95; // @[VTAMemDPI.scala 104:46:@201.10]
  assign _GEN_3 = _T_96 ? 3'h0 : state; // @[VTAMemDPI.scala 104:62:@202.10]
  assign _T_97 = 3'h3 == state; // @[Conditional.scala 37:30:@207.10]
  assign _GEN_4 = io_axi_aw_valid ? 3'h4 : state; // @[VTAMemDPI.scala 109:29:@209.12]
  assign _T_98 = 3'h4 == state; // @[Conditional.scala 37:30:@214.12]
  assign _T_99 = io_axi_w_valid & io_axi_w_bits_last; // @[VTAMemDPI.scala 114:27:@216.14]
  assign _GEN_5 = _T_99 ? 3'h5 : state; // @[VTAMemDPI.scala 114:50:@217.14]
  assign _T_100 = 3'h5 == state; // @[Conditional.scala 37:30:@222.14]
  assign _GEN_6 = io_axi_b_ready ? 3'h0 : state; // @[VTAMemDPI.scala 119:28:@224.16]
  assign _GEN_7 = _T_100 ? _GEN_6 : state; // @[Conditional.scala 39:67:@223.14]
  assign _GEN_8 = _T_98 ? _GEN_5 : _GEN_7; // @[Conditional.scala 39:67:@215.12]
  assign _GEN_9 = _T_97 ? _GEN_4 : _GEN_8; // @[Conditional.scala 39:67:@208.10]
  assign _GEN_10 = _T_92 ? _GEN_3 : _GEN_9; // @[Conditional.scala 39:67:@198.8]
  assign _GEN_11 = _T_91 ? _GEN_2 : _GEN_10; // @[Conditional.scala 39:67:@191.6]
  assign _GEN_12 = _T_90 ? _GEN_1 : _GEN_11; // @[Conditional.scala 40:58:@180.4]
  assign _T_101 = state == 3'h0; // @[VTAMemDPI.scala 125:14:@228.4]
  assign _GEN_13 = io_axi_aw_valid ? 1'h1 : opcode; // @[VTAMemDPI.scala 130:33:@236.8]
  assign _GEN_14 = io_axi_aw_valid ? io_axi_aw_bits_len : len; // @[VTAMemDPI.scala 130:33:@236.8]
  assign _GEN_15 = io_axi_aw_valid ? {{32'd0}, io_axi_aw_bits_addr} : addr; // @[VTAMemDPI.scala 130:33:@236.8]
  assign _GEN_16 = io_axi_ar_valid ? 1'h0 : _GEN_13; // @[VTAMemDPI.scala 126:27:@230.6]
  assign _GEN_17 = io_axi_ar_valid ? io_axi_ar_bits_len : _GEN_14; // @[VTAMemDPI.scala 126:27:@230.6]
  assign _GEN_18 = io_axi_ar_valid ? {{32'd0}, io_axi_ar_bits_addr} : _GEN_15; // @[VTAMemDPI.scala 126:27:@230.6]
  assign _T_104 = state == 3'h2; // @[VTAMemDPI.scala 135:20:@243.6]
  assign _T_107 = len != 8'h0; // @[VTAMemDPI.scala 136:51:@246.8]
  assign _T_108 = _T_93 & _T_107; // @[VTAMemDPI.scala 136:44:@247.8]
  assign _T_110 = len - 8'h1; // @[VTAMemDPI.scala 137:18:@249.10]
  assign _T_111 = $unsigned(_T_110); // @[VTAMemDPI.scala 137:18:@250.10]
  assign _T_112 = _T_111[7:0]; // @[VTAMemDPI.scala 137:18:@251.10]
  assign _GEN_19 = _T_108 ? _T_112 : len; // @[VTAMemDPI.scala 136:60:@248.8]
  assign _GEN_20 = _T_104 ? _GEN_19 : len; // @[VTAMemDPI.scala 135:35:@244.6]
  assign _GEN_21 = _T_101 ? _GEN_16 : opcode; // @[VTAMemDPI.scala 125:25:@229.4]
  assign _GEN_22 = _T_101 ? _GEN_17 : _GEN_20; // @[VTAMemDPI.scala 125:25:@229.4]
  assign _GEN_23 = _T_101 ? _GEN_18 : addr; // @[VTAMemDPI.scala 125:25:@229.4]
  assign _T_113 = state == 3'h1; // @[VTAMemDPI.scala 141:30:@255.4]
  assign _T_114 = _T_113 & io_axi_ar_valid; // @[VTAMemDPI.scala 141:47:@256.4]
  assign _T_115 = state == 3'h3; // @[VTAMemDPI.scala 141:75:@257.4]
  assign _T_116 = _T_115 & io_axi_aw_valid; // @[VTAMemDPI.scala 141:93:@258.4]
  assign _T_129 = state == 3'h4; // @[VTAMemDPI.scala 157:28:@280.4]
  assign io_dpi_req_valid = _T_114 | _T_116; // @[VTAMemDPI.scala 141:20:@260.4]
  assign io_dpi_req_opcode = opcode; // @[VTAMemDPI.scala 142:21:@261.4]
  assign io_dpi_req_len = len; // @[VTAMemDPI.scala 143:18:@262.4]
  assign io_dpi_req_addr = addr; // @[VTAMemDPI.scala 144:19:@263.4]
  assign io_dpi_wr_valid = _T_129 & io_axi_w_valid; // @[VTAMemDPI.scala 157:19:@282.4]
  assign io_dpi_wr_bits = io_axi_w_bits_data; // @[VTAMemDPI.scala 158:18:@283.4]
  assign io_dpi_rd_ready = _T_104 & io_axi_r_ready; // @[VTAMemDPI.scala 155:19:@279.4]
  assign io_axi_aw_ready = state == 3'h3; // @[VTAMemDPI.scala 147:19:@267.4]
  assign io_axi_w_ready = state == 3'h4; // @[VTAMemDPI.scala 159:18:@285.4]
  assign io_axi_b_valid = state == 3'h5; // @[VTAMemDPI.scala 161:18:@287.4]
  assign io_axi_ar_ready = state == 3'h1; // @[VTAMemDPI.scala 146:19:@265.4]
  assign io_axi_r_valid = _T_104 & io_dpi_rd_valid; // @[VTAMemDPI.scala 149:18:@270.4]
  assign io_axi_r_bits_data = io_dpi_rd_bits; // @[VTAMemDPI.scala 150:22:@271.4]
  assign io_axi_r_bits_last = len == 8'h0; // @[VTAMemDPI.scala 151:22:@273.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  opcode = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  len = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  addr = _RAND_2[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      opcode <= 1'h0;
    end else begin
      if (_T_101) begin
        if (io_axi_ar_valid) begin
          opcode <= 1'h0;
        end else begin
          if (io_axi_aw_valid) begin
            opcode <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      len <= 8'h0;
    end else begin
      if (_T_101) begin
        if (io_axi_ar_valid) begin
          len <= io_axi_ar_bits_len;
        end else begin
          if (io_axi_aw_valid) begin
            len <= io_axi_aw_bits_len;
          end
        end
      end else begin
        if (_T_104) begin
          if (_T_108) begin
            len <= _T_112;
          end
        end
      end
    end
    if (reset) begin
      addr <= 64'h0;
    end else begin
      if (_T_101) begin
        if (io_axi_ar_valid) begin
          addr <= {{32'd0}, io_axi_ar_bits_addr};
        end else begin
          if (io_axi_aw_valid) begin
            addr <= {{32'd0}, io_axi_aw_bits_addr};
          end
        end
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_90) begin
        if (io_axi_ar_valid) begin
          state <= 3'h1;
        end else begin
          if (io_axi_aw_valid) begin
            state <= 3'h3;
          end
        end
      end else begin
        if (_T_91) begin
          if (io_axi_ar_valid) begin
            state <= 3'h2;
          end
        end else begin
          if (_T_92) begin
            if (_T_96) begin
              state <= 3'h0;
            end
          end else begin
            if (_T_97) begin
              if (io_axi_aw_valid) begin
                state <= 3'h4;
              end
            end else begin
              if (_T_98) begin
                if (_T_99) begin
                  state <= 3'h5;
                end
              end else begin
                if (_T_100) begin
                  if (io_axi_b_ready) begin
                    state <= 3'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module VTAMem( // @[:@292.2]
  input         clock, // @[:@293.4]
  input         reset, // @[:@294.4]
  output        io_axi_aw_ready, // @[:@295.4]
  input         io_axi_aw_valid, // @[:@295.4]
  input  [31:0] io_axi_aw_bits_addr, // @[:@295.4]
  input  [7:0]  io_axi_aw_bits_len, // @[:@295.4]
  output        io_axi_w_ready, // @[:@295.4]
  input         io_axi_w_valid, // @[:@295.4]
  input  [63:0] io_axi_w_bits_data, // @[:@295.4]
  input         io_axi_w_bits_last, // @[:@295.4]
  input         io_axi_b_ready, // @[:@295.4]
  output        io_axi_b_valid, // @[:@295.4]
  output        io_axi_ar_ready, // @[:@295.4]
  input         io_axi_ar_valid, // @[:@295.4]
  input  [31:0] io_axi_ar_bits_addr, // @[:@295.4]
  input  [7:0]  io_axi_ar_bits_len, // @[:@295.4]
  input         io_axi_r_ready, // @[:@295.4]
  output        io_axi_r_valid, // @[:@295.4]
  output [63:0] io_axi_r_bits_data, // @[:@295.4]
  output        io_axi_r_bits_last // @[:@295.4]
);
  wire  mem_dpi_dpi_req_valid; // @[SimShell.scala 57:23:@297.4]
  wire  mem_dpi_dpi_req_opcode; // @[SimShell.scala 57:23:@297.4]
  wire [7:0] mem_dpi_dpi_req_len; // @[SimShell.scala 57:23:@297.4]
  wire [63:0] mem_dpi_dpi_req_addr; // @[SimShell.scala 57:23:@297.4]
  wire  mem_dpi_dpi_wr_valid; // @[SimShell.scala 57:23:@297.4]
  wire [63:0] mem_dpi_dpi_wr_bits; // @[SimShell.scala 57:23:@297.4]
  wire  mem_dpi_dpi_rd_ready; // @[SimShell.scala 57:23:@297.4]
  wire  mem_dpi_dpi_rd_valid; // @[SimShell.scala 57:23:@297.4]
  wire [63:0] mem_dpi_dpi_rd_bits; // @[SimShell.scala 57:23:@297.4]
  wire  mem_dpi_reset; // @[SimShell.scala 57:23:@297.4]
  wire  mem_dpi_clock; // @[SimShell.scala 57:23:@297.4]
  wire  mem_axi_clock; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_reset; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_dpi_req_valid; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_dpi_req_opcode; // @[SimShell.scala 58:23:@301.4]
  wire [7:0] mem_axi_io_dpi_req_len; // @[SimShell.scala 58:23:@301.4]
  wire [63:0] mem_axi_io_dpi_req_addr; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_dpi_wr_valid; // @[SimShell.scala 58:23:@301.4]
  wire [63:0] mem_axi_io_dpi_wr_bits; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_dpi_rd_ready; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_dpi_rd_valid; // @[SimShell.scala 58:23:@301.4]
  wire [63:0] mem_axi_io_dpi_rd_bits; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_aw_ready; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_aw_valid; // @[SimShell.scala 58:23:@301.4]
  wire [31:0] mem_axi_io_axi_aw_bits_addr; // @[SimShell.scala 58:23:@301.4]
  wire [7:0] mem_axi_io_axi_aw_bits_len; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_w_ready; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_w_valid; // @[SimShell.scala 58:23:@301.4]
  wire [63:0] mem_axi_io_axi_w_bits_data; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_w_bits_last; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_b_ready; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_b_valid; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_ar_ready; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_ar_valid; // @[SimShell.scala 58:23:@301.4]
  wire [31:0] mem_axi_io_axi_ar_bits_addr; // @[SimShell.scala 58:23:@301.4]
  wire [7:0] mem_axi_io_axi_ar_bits_len; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_r_ready; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_r_valid; // @[SimShell.scala 58:23:@301.4]
  wire [63:0] mem_axi_io_axi_r_bits_data; // @[SimShell.scala 58:23:@301.4]
  wire  mem_axi_io_axi_r_bits_last; // @[SimShell.scala 58:23:@301.4]
  VTAMemDPI mem_dpi ( // @[SimShell.scala 57:23:@297.4]
    .dpi_req_valid(mem_dpi_dpi_req_valid),
    .dpi_req_opcode(mem_dpi_dpi_req_opcode),
    .dpi_req_len(mem_dpi_dpi_req_len),
    .dpi_req_addr(mem_dpi_dpi_req_addr),
    .dpi_wr_valid(mem_dpi_dpi_wr_valid),
    .dpi_wr_bits(mem_dpi_dpi_wr_bits),
    .dpi_rd_ready(mem_dpi_dpi_rd_ready),
    .dpi_rd_valid(mem_dpi_dpi_rd_valid),
    .dpi_rd_bits(mem_dpi_dpi_rd_bits),
    .reset(mem_dpi_reset),
    .clock(mem_dpi_clock)
  );
  VTAMemDPIToAXI mem_axi ( // @[SimShell.scala 58:23:@301.4]
    .clock(mem_axi_clock),
    .reset(mem_axi_reset),
    .io_dpi_req_valid(mem_axi_io_dpi_req_valid),
    .io_dpi_req_opcode(mem_axi_io_dpi_req_opcode),
    .io_dpi_req_len(mem_axi_io_dpi_req_len),
    .io_dpi_req_addr(mem_axi_io_dpi_req_addr),
    .io_dpi_wr_valid(mem_axi_io_dpi_wr_valid),
    .io_dpi_wr_bits(mem_axi_io_dpi_wr_bits),
    .io_dpi_rd_ready(mem_axi_io_dpi_rd_ready),
    .io_dpi_rd_valid(mem_axi_io_dpi_rd_valid),
    .io_dpi_rd_bits(mem_axi_io_dpi_rd_bits),
    .io_axi_aw_ready(mem_axi_io_axi_aw_ready),
    .io_axi_aw_valid(mem_axi_io_axi_aw_valid),
    .io_axi_aw_bits_addr(mem_axi_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(mem_axi_io_axi_aw_bits_len),
    .io_axi_w_ready(mem_axi_io_axi_w_ready),
    .io_axi_w_valid(mem_axi_io_axi_w_valid),
    .io_axi_w_bits_data(mem_axi_io_axi_w_bits_data),
    .io_axi_w_bits_last(mem_axi_io_axi_w_bits_last),
    .io_axi_b_ready(mem_axi_io_axi_b_ready),
    .io_axi_b_valid(mem_axi_io_axi_b_valid),
    .io_axi_ar_ready(mem_axi_io_axi_ar_ready),
    .io_axi_ar_valid(mem_axi_io_axi_ar_valid),
    .io_axi_ar_bits_addr(mem_axi_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(mem_axi_io_axi_ar_bits_len),
    .io_axi_r_ready(mem_axi_io_axi_r_ready),
    .io_axi_r_valid(mem_axi_io_axi_r_valid),
    .io_axi_r_bits_data(mem_axi_io_axi_r_bits_data),
    .io_axi_r_bits_last(mem_axi_io_axi_r_bits_last)
  );
  assign io_axi_aw_ready = mem_axi_io_axi_aw_ready; // @[SimShell.scala 62:18:@359.4]
  assign io_axi_w_ready = mem_axi_io_axi_w_ready; // @[SimShell.scala 62:18:@346.4]
  assign io_axi_b_valid = mem_axi_io_axi_b_valid; // @[SimShell.scala 62:18:@338.4]
  assign io_axi_ar_ready = mem_axi_io_axi_ar_ready; // @[SimShell.scala 62:18:@334.4]
  assign io_axi_r_valid = mem_axi_io_axi_r_valid; // @[SimShell.scala 62:18:@320.4]
  assign io_axi_r_bits_data = mem_axi_io_axi_r_bits_data; // @[SimShell.scala 62:18:@319.4]
  assign io_axi_r_bits_last = mem_axi_io_axi_r_bits_last; // @[SimShell.scala 62:18:@317.4]
  assign mem_dpi_dpi_req_valid = mem_axi_io_dpi_req_valid; // @[SimShell.scala 61:18:@314.4]
  assign mem_dpi_dpi_req_opcode = mem_axi_io_dpi_req_opcode; // @[SimShell.scala 61:18:@313.4]
  assign mem_dpi_dpi_req_len = mem_axi_io_dpi_req_len; // @[SimShell.scala 61:18:@312.4]
  assign mem_dpi_dpi_req_addr = mem_axi_io_dpi_req_addr; // @[SimShell.scala 61:18:@311.4]
  assign mem_dpi_dpi_wr_valid = mem_axi_io_dpi_wr_valid; // @[SimShell.scala 61:18:@310.4]
  assign mem_dpi_dpi_wr_bits = mem_axi_io_dpi_wr_bits; // @[SimShell.scala 61:18:@309.4]
  assign mem_dpi_dpi_rd_ready = mem_axi_io_dpi_rd_ready; // @[SimShell.scala 61:18:@308.4]
  assign mem_dpi_reset = reset; // @[SimShell.scala 59:20:@304.4]
  assign mem_dpi_clock = clock; // @[SimShell.scala 60:20:@305.4]
  assign mem_axi_clock = clock; // @[:@302.4]
  assign mem_axi_reset = reset; // @[:@303.4]
  assign mem_axi_io_dpi_rd_valid = mem_dpi_dpi_rd_valid; // @[SimShell.scala 61:18:@307.4]
  assign mem_axi_io_dpi_rd_bits = mem_dpi_dpi_rd_bits; // @[SimShell.scala 61:18:@306.4]
  assign mem_axi_io_axi_aw_valid = io_axi_aw_valid; // @[SimShell.scala 62:18:@358.4]
  assign mem_axi_io_axi_aw_bits_addr = io_axi_aw_bits_addr; // @[SimShell.scala 62:18:@357.4]
  assign mem_axi_io_axi_aw_bits_len = io_axi_aw_bits_len; // @[SimShell.scala 62:18:@354.4]
  assign mem_axi_io_axi_w_valid = io_axi_w_valid; // @[SimShell.scala 62:18:@345.4]
  assign mem_axi_io_axi_w_bits_data = io_axi_w_bits_data; // @[SimShell.scala 62:18:@344.4]
  assign mem_axi_io_axi_w_bits_last = io_axi_w_bits_last; // @[SimShell.scala 62:18:@342.4]
  assign mem_axi_io_axi_b_ready = io_axi_b_ready; // @[SimShell.scala 62:18:@339.4]
  assign mem_axi_io_axi_ar_valid = io_axi_ar_valid; // @[SimShell.scala 62:18:@333.4]
  assign mem_axi_io_axi_ar_bits_addr = io_axi_ar_bits_addr; // @[SimShell.scala 62:18:@332.4]
  assign mem_axi_io_axi_ar_bits_len = io_axi_ar_bits_len; // @[SimShell.scala 62:18:@329.4]
  assign mem_axi_io_axi_r_ready = io_axi_r_ready; // @[SimShell.scala 62:18:@321.4]
endmodule
module SimShell( // @[:@361.2]
  input         clock, // @[:@362.4]
  input         reset, // @[:@363.4]
  output        mem_aw_ready, // @[:@364.4]
  input         mem_aw_valid, // @[:@364.4]
  input  [31:0] mem_aw_bits_addr, // @[:@364.4]
  input  [7:0]  mem_aw_bits_len, // @[:@364.4]
  output        mem_w_ready, // @[:@364.4]
  input         mem_w_valid, // @[:@364.4]
  input  [63:0] mem_w_bits_data, // @[:@364.4]
  input         mem_w_bits_last, // @[:@364.4]
  input         mem_b_ready, // @[:@364.4]
  output        mem_b_valid, // @[:@364.4]
  output        mem_ar_ready, // @[:@364.4]
  input         mem_ar_valid, // @[:@364.4]
  input  [31:0] mem_ar_bits_addr, // @[:@364.4]
  input  [7:0]  mem_ar_bits_len, // @[:@364.4]
  input         mem_r_ready, // @[:@364.4]
  output        mem_r_valid, // @[:@364.4]
  output [63:0] mem_r_bits_data, // @[:@364.4]
  output        mem_r_bits_last, // @[:@364.4]
  input         host_aw_ready, // @[:@365.4]
  output        host_aw_valid, // @[:@365.4]
  output [15:0] host_aw_bits_addr, // @[:@365.4]
  input         host_w_ready, // @[:@365.4]
  output        host_w_valid, // @[:@365.4]
  output [31:0] host_w_bits_data, // @[:@365.4]
  output        host_b_ready, // @[:@365.4]
  input         host_b_valid, // @[:@365.4]
  input         host_ar_ready, // @[:@365.4]
  output        host_ar_valid, // @[:@365.4]
  output [15:0] host_ar_bits_addr, // @[:@365.4]
  output        host_r_ready, // @[:@365.4]
  input         host_r_valid, // @[:@365.4]
  input  [31:0] host_r_bits_data, // @[:@365.4]
  input         sim_clock, // @[:@366.4]
  output        sim_wait // @[:@367.4]
);
  wire  mod_sim_clock; // @[SimShell.scala 91:23:@369.4]
  wire  mod_sim_reset; // @[SimShell.scala 91:23:@369.4]
  wire  mod_sim_sim_wait; // @[SimShell.scala 91:23:@369.4]
  wire  mod_host_clock; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_reset; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_aw_ready; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_aw_valid; // @[SimShell.scala 92:24:@372.4]
  wire [15:0] mod_host_io_axi_aw_bits_addr; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_w_ready; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_w_valid; // @[SimShell.scala 92:24:@372.4]
  wire [31:0] mod_host_io_axi_w_bits_data; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_b_ready; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_b_valid; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_ar_ready; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_ar_valid; // @[SimShell.scala 92:24:@372.4]
  wire [15:0] mod_host_io_axi_ar_bits_addr; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_r_ready; // @[SimShell.scala 92:24:@372.4]
  wire  mod_host_io_axi_r_valid; // @[SimShell.scala 92:24:@372.4]
  wire [31:0] mod_host_io_axi_r_bits_data; // @[SimShell.scala 92:24:@372.4]
  wire  mod_mem_clock; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_reset; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_aw_ready; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_aw_valid; // @[SimShell.scala 93:23:@375.4]
  wire [31:0] mod_mem_io_axi_aw_bits_addr; // @[SimShell.scala 93:23:@375.4]
  wire [7:0] mod_mem_io_axi_aw_bits_len; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_w_ready; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_w_valid; // @[SimShell.scala 93:23:@375.4]
  wire [63:0] mod_mem_io_axi_w_bits_data; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_w_bits_last; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_b_ready; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_b_valid; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_ar_ready; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_ar_valid; // @[SimShell.scala 93:23:@375.4]
  wire [31:0] mod_mem_io_axi_ar_bits_addr; // @[SimShell.scala 93:23:@375.4]
  wire [7:0] mod_mem_io_axi_ar_bits_len; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_r_ready; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_r_valid; // @[SimShell.scala 93:23:@375.4]
  wire [63:0] mod_mem_io_axi_r_bits_data; // @[SimShell.scala 93:23:@375.4]
  wire  mod_mem_io_axi_r_bits_last; // @[SimShell.scala 93:23:@375.4]
  VTASim mod_sim ( // @[SimShell.scala 91:23:@369.4]
    .clock(mod_sim_clock),
    .reset(mod_sim_reset),
    .sim_wait(mod_sim_sim_wait)
  );
  VTAHost mod_host ( // @[SimShell.scala 92:24:@372.4]
    .clock(mod_host_clock),
    .reset(mod_host_reset),
    .io_axi_aw_ready(mod_host_io_axi_aw_ready),
    .io_axi_aw_valid(mod_host_io_axi_aw_valid),
    .io_axi_aw_bits_addr(mod_host_io_axi_aw_bits_addr),
    .io_axi_w_ready(mod_host_io_axi_w_ready),
    .io_axi_w_valid(mod_host_io_axi_w_valid),
    .io_axi_w_bits_data(mod_host_io_axi_w_bits_data),
    .io_axi_b_ready(mod_host_io_axi_b_ready),
    .io_axi_b_valid(mod_host_io_axi_b_valid),
    .io_axi_ar_ready(mod_host_io_axi_ar_ready),
    .io_axi_ar_valid(mod_host_io_axi_ar_valid),
    .io_axi_ar_bits_addr(mod_host_io_axi_ar_bits_addr),
    .io_axi_r_ready(mod_host_io_axi_r_ready),
    .io_axi_r_valid(mod_host_io_axi_r_valid),
    .io_axi_r_bits_data(mod_host_io_axi_r_bits_data)
  );
  VTAMem mod_mem ( // @[SimShell.scala 93:23:@375.4]
    .clock(mod_mem_clock),
    .reset(mod_mem_reset),
    .io_axi_aw_ready(mod_mem_io_axi_aw_ready),
    .io_axi_aw_valid(mod_mem_io_axi_aw_valid),
    .io_axi_aw_bits_addr(mod_mem_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(mod_mem_io_axi_aw_bits_len),
    .io_axi_w_ready(mod_mem_io_axi_w_ready),
    .io_axi_w_valid(mod_mem_io_axi_w_valid),
    .io_axi_w_bits_data(mod_mem_io_axi_w_bits_data),
    .io_axi_w_bits_last(mod_mem_io_axi_w_bits_last),
    .io_axi_b_ready(mod_mem_io_axi_b_ready),
    .io_axi_b_valid(mod_mem_io_axi_b_valid),
    .io_axi_ar_ready(mod_mem_io_axi_ar_ready),
    .io_axi_ar_valid(mod_mem_io_axi_ar_valid),
    .io_axi_ar_bits_addr(mod_mem_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(mod_mem_io_axi_ar_bits_len),
    .io_axi_r_ready(mod_mem_io_axi_r_ready),
    .io_axi_r_valid(mod_mem_io_axi_r_valid),
    .io_axi_r_bits_data(mod_mem_io_axi_r_bits_data),
    .io_axi_r_bits_last(mod_mem_io_axi_r_bits_last)
  );
  assign mem_aw_ready = mod_mem_io_axi_aw_ready; // @[SimShell.scala 94:7:@422.4]
  assign mem_w_ready = mod_mem_io_axi_w_ready; // @[SimShell.scala 94:7:@409.4]
  assign mem_b_valid = mod_mem_io_axi_b_valid; // @[SimShell.scala 94:7:@401.4]
  assign mem_ar_ready = mod_mem_io_axi_ar_ready; // @[SimShell.scala 94:7:@397.4]
  assign mem_r_valid = mod_mem_io_axi_r_valid; // @[SimShell.scala 94:7:@383.4]
  assign mem_r_bits_data = mod_mem_io_axi_r_bits_data; // @[SimShell.scala 94:7:@382.4]
  assign mem_r_bits_last = mod_mem_io_axi_r_bits_last; // @[SimShell.scala 94:7:@380.4]
  assign host_aw_valid = mod_host_io_axi_aw_valid; // @[SimShell.scala 95:8:@438.4]
  assign host_aw_bits_addr = mod_host_io_axi_aw_bits_addr; // @[SimShell.scala 95:8:@437.4]
  assign host_w_valid = mod_host_io_axi_w_valid; // @[SimShell.scala 95:8:@435.4]
  assign host_w_bits_data = mod_host_io_axi_w_bits_data; // @[SimShell.scala 95:8:@434.4]
  assign host_b_ready = mod_host_io_axi_b_ready; // @[SimShell.scala 95:8:@432.4]
  assign host_ar_valid = mod_host_io_axi_ar_valid; // @[SimShell.scala 95:8:@428.4]
  assign host_ar_bits_addr = mod_host_io_axi_ar_bits_addr; // @[SimShell.scala 95:8:@427.4]
  assign host_r_ready = mod_host_io_axi_r_ready; // @[SimShell.scala 95:8:@426.4]
  assign sim_wait = mod_sim_sim_wait; // @[SimShell.scala 98:12:@442.4]
  assign mod_sim_clock = sim_clock; // @[:@370.4 SimShell.scala 97:17:@441.4]
  assign mod_sim_reset = reset; // @[:@371.4 SimShell.scala 96:17:@440.4]
  assign mod_host_clock = clock; // @[:@373.4]
  assign mod_host_reset = reset; // @[:@374.4]
  assign mod_host_io_axi_aw_ready = host_aw_ready; // @[SimShell.scala 95:8:@439.4]
  assign mod_host_io_axi_w_ready = host_w_ready; // @[SimShell.scala 95:8:@436.4]
  assign mod_host_io_axi_b_valid = host_b_valid; // @[SimShell.scala 95:8:@431.4]
  assign mod_host_io_axi_ar_ready = host_ar_ready; // @[SimShell.scala 95:8:@429.4]
  assign mod_host_io_axi_r_valid = host_r_valid; // @[SimShell.scala 95:8:@425.4]
  assign mod_host_io_axi_r_bits_data = host_r_bits_data; // @[SimShell.scala 95:8:@424.4]
  assign mod_mem_clock = clock; // @[:@376.4]
  assign mod_mem_reset = reset; // @[:@377.4]
  assign mod_mem_io_axi_aw_valid = mem_aw_valid; // @[SimShell.scala 94:7:@421.4]
  assign mod_mem_io_axi_aw_bits_addr = mem_aw_bits_addr; // @[SimShell.scala 94:7:@420.4]
  assign mod_mem_io_axi_aw_bits_len = mem_aw_bits_len; // @[SimShell.scala 94:7:@417.4]
  assign mod_mem_io_axi_w_valid = mem_w_valid; // @[SimShell.scala 94:7:@408.4]
  assign mod_mem_io_axi_w_bits_data = mem_w_bits_data; // @[SimShell.scala 94:7:@407.4]
  assign mod_mem_io_axi_w_bits_last = mem_w_bits_last; // @[SimShell.scala 94:7:@405.4]
  assign mod_mem_io_axi_b_ready = mem_b_ready; // @[SimShell.scala 94:7:@402.4]
  assign mod_mem_io_axi_ar_valid = mem_ar_valid; // @[SimShell.scala 94:7:@396.4]
  assign mod_mem_io_axi_ar_bits_addr = mem_ar_bits_addr; // @[SimShell.scala 94:7:@395.4]
  assign mod_mem_io_axi_ar_bits_len = mem_ar_bits_len; // @[SimShell.scala 94:7:@392.4]
  assign mod_mem_io_axi_r_ready = mem_r_ready; // @[SimShell.scala 94:7:@384.4]
endmodule
module VCR( // @[:@444.2]
  input         clock, // @[:@445.4]
  input         reset, // @[:@446.4]
  output        io_host_aw_ready, // @[:@447.4]
  input         io_host_aw_valid, // @[:@447.4]
  input  [15:0] io_host_aw_bits_addr, // @[:@447.4]
  output        io_host_w_ready, // @[:@447.4]
  input         io_host_w_valid, // @[:@447.4]
  input  [31:0] io_host_w_bits_data, // @[:@447.4]
  input         io_host_b_ready, // @[:@447.4]
  output        io_host_b_valid, // @[:@447.4]
  output        io_host_ar_ready, // @[:@447.4]
  input         io_host_ar_valid, // @[:@447.4]
  input  [15:0] io_host_ar_bits_addr, // @[:@447.4]
  input         io_host_r_ready, // @[:@447.4]
  output        io_host_r_valid, // @[:@447.4]
  output [31:0] io_host_r_bits_data, // @[:@447.4]
  output        io_vcr_launch, // @[:@447.4]
  input         io_vcr_finish, // @[:@447.4]
  input         io_vcr_ecnt_0_valid, // @[:@447.4]
  input  [31:0] io_vcr_ecnt_0_bits, // @[:@447.4]
  output [31:0] io_vcr_vals_0, // @[:@447.4]
  output [31:0] io_vcr_ptrs_0, // @[:@447.4]
  output [31:0] io_vcr_ptrs_1, // @[:@447.4]
  output [31:0] io_vcr_ptrs_2, // @[:@447.4]
  output [31:0] io_vcr_ptrs_3, // @[:@447.4]
  output [31:0] io_vcr_ptrs_4, // @[:@447.4]
  output [31:0] io_vcr_ptrs_5, // @[:@447.4]
  input         io_vcr_ucnt_0_valid, // @[:@447.4]
  input  [31:0] io_vcr_ucnt_0_bits // @[:@447.4]
);
  reg [15:0] waddr; // @[VCR.scala 94:22:@449.4]
  reg [31:0] _RAND_0;
  reg [1:0] wstate; // @[VCR.scala 97:23:@450.4]
  reg [31:0] _RAND_1;
  reg  rstate; // @[VCR.scala 101:23:@451.4]
  reg [31:0] _RAND_2;
  reg [31:0] rdata; // @[VCR.scala 102:22:@452.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_0; // @[VCR.scala 108:37:@453.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_1; // @[VCR.scala 108:37:@454.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_2; // @[VCR.scala 108:37:@455.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_3; // @[VCR.scala 108:37:@456.4]
  reg [31:0] _RAND_7;
  reg [31:0] reg_4; // @[VCR.scala 108:37:@457.4]
  reg [31:0] _RAND_8;
  reg [31:0] reg_5; // @[VCR.scala 108:37:@458.4]
  reg [31:0] _RAND_9;
  reg [31:0] reg_6; // @[VCR.scala 108:37:@459.4]
  reg [31:0] _RAND_10;
  reg [31:0] reg_7; // @[VCR.scala 108:37:@460.4]
  reg [31:0] _RAND_11;
  reg [31:0] reg_8; // @[VCR.scala 108:37:@461.4]
  reg [31:0] _RAND_12;
  reg [31:0] reg_9; // @[VCR.scala 108:37:@462.4]
  reg [31:0] _RAND_13;
  wire  _T_159; // @[Conditional.scala 37:30:@463.4]
  wire [1:0] _GEN_0; // @[VCR.scala 118:30:@465.6]
  wire  _T_160; // @[Conditional.scala 37:30:@470.6]
  wire [1:0] _GEN_1; // @[VCR.scala 123:29:@472.8]
  wire  _T_161; // @[Conditional.scala 37:30:@477.8]
  wire [1:0] _GEN_2; // @[VCR.scala 128:29:@479.10]
  wire [1:0] _GEN_3; // @[Conditional.scala 39:67:@478.8]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@471.6]
  wire [1:0] _GEN_5; // @[Conditional.scala 40:58:@464.4]
  wire  _T_162; // @[Decoupled.scala 37:37:@483.4]
  wire [15:0] _GEN_6; // @[VCR.scala 134:27:@484.4]
  wire  _T_167; // @[Conditional.scala 37:30:@494.4]
  wire  _GEN_7; // @[VCR.scala 143:30:@496.6]
  wire  _GEN_8; // @[VCR.scala 148:29:@503.8]
  wire  _GEN_9; // @[Conditional.scala 39:67:@502.6]
  wire  _GEN_10; // @[Conditional.scala 40:58:@495.4]
  wire  _T_173; // @[Decoupled.scala 37:37:@517.6]
  wire  _T_175; // @[VCR.scala 161:44:@518.6]
  wire  _T_176; // @[VCR.scala 161:31:@519.6]
  wire [31:0] _GEN_11; // @[VCR.scala 161:55:@520.6]
  wire [31:0] _GEN_12; // @[VCR.scala 159:23:@513.4]
  wire  _T_179; // @[VCR.scala 168:51:@528.6]
  wire  _T_180; // @[VCR.scala 168:33:@529.6]
  wire [31:0] _GEN_13; // @[VCR.scala 168:62:@530.6]
  wire [31:0] _GEN_14; // @[VCR.scala 166:32:@523.4]
  wire  _T_183; // @[VCR.scala 174:45:@534.4]
  wire  _T_184; // @[VCR.scala 174:27:@535.4]
  wire [31:0] _GEN_15; // @[VCR.scala 174:56:@536.4]
  wire  _T_187; // @[VCR.scala 174:45:@540.4]
  wire  _T_188; // @[VCR.scala 174:27:@541.4]
  wire [31:0] _GEN_16; // @[VCR.scala 174:56:@542.4]
  wire  _T_191; // @[VCR.scala 174:45:@546.4]
  wire  _T_192; // @[VCR.scala 174:27:@547.4]
  wire [31:0] _GEN_17; // @[VCR.scala 174:56:@548.4]
  wire  _T_195; // @[VCR.scala 174:45:@552.4]
  wire  _T_196; // @[VCR.scala 174:27:@553.4]
  wire [31:0] _GEN_18; // @[VCR.scala 174:56:@554.4]
  wire  _T_199; // @[VCR.scala 174:45:@558.4]
  wire  _T_200; // @[VCR.scala 174:27:@559.4]
  wire [31:0] _GEN_19; // @[VCR.scala 174:56:@560.4]
  wire  _T_203; // @[VCR.scala 174:45:@564.4]
  wire  _T_204; // @[VCR.scala 174:27:@565.4]
  wire [31:0] _GEN_20; // @[VCR.scala 174:56:@566.4]
  wire  _T_207; // @[VCR.scala 174:45:@570.4]
  wire  _T_208; // @[VCR.scala 174:27:@571.4]
  wire [31:0] _GEN_21; // @[VCR.scala 174:56:@572.4]
  wire  _T_209; // @[Decoupled.scala 37:37:@575.4]
  wire  _T_211; // @[Mux.scala 46:19:@577.6]
  wire [31:0] _T_212; // @[Mux.scala 46:16:@578.6]
  wire  _T_213; // @[Mux.scala 46:19:@579.6]
  wire [31:0] _T_214; // @[Mux.scala 46:16:@580.6]
  wire  _T_215; // @[Mux.scala 46:19:@581.6]
  wire [31:0] _T_216; // @[Mux.scala 46:16:@582.6]
  wire  _T_217; // @[Mux.scala 46:19:@583.6]
  wire [31:0] _T_218; // @[Mux.scala 46:16:@584.6]
  wire  _T_219; // @[Mux.scala 46:19:@585.6]
  wire [31:0] _T_220; // @[Mux.scala 46:16:@586.6]
  wire  _T_221; // @[Mux.scala 46:19:@587.6]
  wire [31:0] _T_222; // @[Mux.scala 46:16:@588.6]
  wire  _T_223; // @[Mux.scala 46:19:@589.6]
  wire [31:0] _T_224; // @[Mux.scala 46:16:@590.6]
  wire  _T_225; // @[Mux.scala 46:19:@591.6]
  wire [31:0] _T_226; // @[Mux.scala 46:16:@592.6]
  wire  _T_227; // @[Mux.scala 46:19:@593.6]
  wire [31:0] _T_228; // @[Mux.scala 46:16:@594.6]
  wire  _T_229; // @[Mux.scala 46:19:@595.6]
  wire [31:0] _T_230; // @[Mux.scala 46:16:@596.6]
  wire [31:0] _GEN_22; // @[VCR.scala 179:27:@576.4]
  wire  _T_234; // @[VCR.scala 202:51:@613.6]
  wire  _T_235; // @[VCR.scala 202:33:@614.6]
  wire [31:0] _GEN_23; // @[VCR.scala 202:62:@615.6]
  wire [31:0] _GEN_24; // @[VCR.scala 200:32:@608.4]
  assign _T_159 = 2'h0 == wstate; // @[Conditional.scala 37:30:@463.4]
  assign _GEN_0 = io_host_aw_valid ? 2'h1 : wstate; // @[VCR.scala 118:30:@465.6]
  assign _T_160 = 2'h1 == wstate; // @[Conditional.scala 37:30:@470.6]
  assign _GEN_1 = io_host_w_valid ? 2'h2 : wstate; // @[VCR.scala 123:29:@472.8]
  assign _T_161 = 2'h2 == wstate; // @[Conditional.scala 37:30:@477.8]
  assign _GEN_2 = io_host_b_ready ? 2'h0 : wstate; // @[VCR.scala 128:29:@479.10]
  assign _GEN_3 = _T_161 ? _GEN_2 : wstate; // @[Conditional.scala 39:67:@478.8]
  assign _GEN_4 = _T_160 ? _GEN_1 : _GEN_3; // @[Conditional.scala 39:67:@471.6]
  assign _GEN_5 = _T_159 ? _GEN_0 : _GEN_4; // @[Conditional.scala 40:58:@464.4]
  assign _T_162 = io_host_aw_ready & io_host_aw_valid; // @[Decoupled.scala 37:37:@483.4]
  assign _GEN_6 = _T_162 ? io_host_aw_bits_addr : waddr; // @[VCR.scala 134:27:@484.4]
  assign _T_167 = 1'h0 == rstate; // @[Conditional.scala 37:30:@494.4]
  assign _GEN_7 = io_host_ar_valid ? 1'h1 : rstate; // @[VCR.scala 143:30:@496.6]
  assign _GEN_8 = io_host_r_ready ? 1'h0 : rstate; // @[VCR.scala 148:29:@503.8]
  assign _GEN_9 = rstate ? _GEN_8 : rstate; // @[Conditional.scala 39:67:@502.6]
  assign _GEN_10 = _T_167 ? _GEN_7 : _GEN_9; // @[Conditional.scala 40:58:@495.4]
  assign _T_173 = io_host_w_ready & io_host_w_valid; // @[Decoupled.scala 37:37:@517.6]
  assign _T_175 = 16'h0 == waddr; // @[VCR.scala 161:44:@518.6]
  assign _T_176 = _T_173 & _T_175; // @[VCR.scala 161:31:@519.6]
  assign _GEN_11 = _T_176 ? io_host_w_bits_data : reg_0; // @[VCR.scala 161:55:@520.6]
  assign _GEN_12 = io_vcr_finish ? 32'h2 : _GEN_11; // @[VCR.scala 159:23:@513.4]
  assign _T_179 = 16'h4 == waddr; // @[VCR.scala 168:51:@528.6]
  assign _T_180 = _T_173 & _T_179; // @[VCR.scala 168:33:@529.6]
  assign _GEN_13 = _T_180 ? io_host_w_bits_data : reg_1; // @[VCR.scala 168:62:@530.6]
  assign _GEN_14 = io_vcr_ecnt_0_valid ? io_vcr_ecnt_0_bits : _GEN_13; // @[VCR.scala 166:32:@523.4]
  assign _T_183 = 16'h8 == waddr; // @[VCR.scala 174:45:@534.4]
  assign _T_184 = _T_173 & _T_183; // @[VCR.scala 174:27:@535.4]
  assign _GEN_15 = _T_184 ? io_host_w_bits_data : reg_2; // @[VCR.scala 174:56:@536.4]
  assign _T_187 = 16'hc == waddr; // @[VCR.scala 174:45:@540.4]
  assign _T_188 = _T_173 & _T_187; // @[VCR.scala 174:27:@541.4]
  assign _GEN_16 = _T_188 ? io_host_w_bits_data : reg_3; // @[VCR.scala 174:56:@542.4]
  assign _T_191 = 16'h10 == waddr; // @[VCR.scala 174:45:@546.4]
  assign _T_192 = _T_173 & _T_191; // @[VCR.scala 174:27:@547.4]
  assign _GEN_17 = _T_192 ? io_host_w_bits_data : reg_4; // @[VCR.scala 174:56:@548.4]
  assign _T_195 = 16'h14 == waddr; // @[VCR.scala 174:45:@552.4]
  assign _T_196 = _T_173 & _T_195; // @[VCR.scala 174:27:@553.4]
  assign _GEN_18 = _T_196 ? io_host_w_bits_data : reg_5; // @[VCR.scala 174:56:@554.4]
  assign _T_199 = 16'h18 == waddr; // @[VCR.scala 174:45:@558.4]
  assign _T_200 = _T_173 & _T_199; // @[VCR.scala 174:27:@559.4]
  assign _GEN_19 = _T_200 ? io_host_w_bits_data : reg_6; // @[VCR.scala 174:56:@560.4]
  assign _T_203 = 16'h1c == waddr; // @[VCR.scala 174:45:@564.4]
  assign _T_204 = _T_173 & _T_203; // @[VCR.scala 174:27:@565.4]
  assign _GEN_20 = _T_204 ? io_host_w_bits_data : reg_7; // @[VCR.scala 174:56:@566.4]
  assign _T_207 = 16'h20 == waddr; // @[VCR.scala 174:45:@570.4]
  assign _T_208 = _T_173 & _T_207; // @[VCR.scala 174:27:@571.4]
  assign _GEN_21 = _T_208 ? io_host_w_bits_data : reg_8; // @[VCR.scala 174:56:@572.4]
  assign _T_209 = io_host_ar_ready & io_host_ar_valid; // @[Decoupled.scala 37:37:@575.4]
  assign _T_211 = 16'h24 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@577.6]
  assign _T_212 = _T_211 ? reg_9 : 32'h0; // @[Mux.scala 46:16:@578.6]
  assign _T_213 = 16'h20 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@579.6]
  assign _T_214 = _T_213 ? reg_8 : _T_212; // @[Mux.scala 46:16:@580.6]
  assign _T_215 = 16'h1c == io_host_ar_bits_addr; // @[Mux.scala 46:19:@581.6]
  assign _T_216 = _T_215 ? reg_7 : _T_214; // @[Mux.scala 46:16:@582.6]
  assign _T_217 = 16'h18 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@583.6]
  assign _T_218 = _T_217 ? reg_6 : _T_216; // @[Mux.scala 46:16:@584.6]
  assign _T_219 = 16'h14 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@585.6]
  assign _T_220 = _T_219 ? reg_5 : _T_218; // @[Mux.scala 46:16:@586.6]
  assign _T_221 = 16'h10 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@587.6]
  assign _T_222 = _T_221 ? reg_4 : _T_220; // @[Mux.scala 46:16:@588.6]
  assign _T_223 = 16'hc == io_host_ar_bits_addr; // @[Mux.scala 46:19:@589.6]
  assign _T_224 = _T_223 ? reg_3 : _T_222; // @[Mux.scala 46:16:@590.6]
  assign _T_225 = 16'h8 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@591.6]
  assign _T_226 = _T_225 ? reg_2 : _T_224; // @[Mux.scala 46:16:@592.6]
  assign _T_227 = 16'h4 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@593.6]
  assign _T_228 = _T_227 ? reg_1 : _T_226; // @[Mux.scala 46:16:@594.6]
  assign _T_229 = 16'h0 == io_host_ar_bits_addr; // @[Mux.scala 46:19:@595.6]
  assign _T_230 = _T_229 ? reg_0 : _T_228; // @[Mux.scala 46:16:@596.6]
  assign _GEN_22 = _T_209 ? _T_230 : rdata; // @[VCR.scala 179:27:@576.4]
  assign _T_234 = 16'h24 == waddr; // @[VCR.scala 202:51:@613.6]
  assign _T_235 = _T_173 & _T_234; // @[VCR.scala 202:33:@614.6]
  assign _GEN_23 = _T_235 ? io_host_w_bits_data : reg_9; // @[VCR.scala 202:62:@615.6]
  assign _GEN_24 = io_vcr_ucnt_0_valid ? io_vcr_ucnt_0_bits : _GEN_23; // @[VCR.scala 200:32:@608.4]
  assign io_host_aw_ready = wstate == 2'h0; // @[VCR.scala 136:20:@488.4]
  assign io_host_w_ready = wstate == 2'h1; // @[VCR.scala 137:19:@490.4]
  assign io_host_b_valid = wstate == 2'h2; // @[VCR.scala 138:19:@492.4]
  assign io_host_ar_ready = rstate == 1'h0; // @[VCR.scala 154:20:@508.4]
  assign io_host_r_valid = rstate; // @[VCR.scala 155:19:@510.4]
  assign io_host_r_bits_data = rdata; // @[VCR.scala 156:23:@511.4]
  assign io_vcr_launch = reg_0[0]; // @[VCR.scala 183:17:@600.4]
  assign io_vcr_vals_0 = reg_2; // @[VCR.scala 186:20:@601.4]
  assign io_vcr_ptrs_0 = reg_3; // @[VCR.scala 191:22:@602.4]
  assign io_vcr_ptrs_1 = reg_4; // @[VCR.scala 191:22:@603.4]
  assign io_vcr_ptrs_2 = reg_5; // @[VCR.scala 191:22:@604.4]
  assign io_vcr_ptrs_3 = reg_6; // @[VCR.scala 191:22:@605.4]
  assign io_vcr_ptrs_4 = reg_7; // @[VCR.scala 191:22:@606.4]
  assign io_vcr_ptrs_5 = reg_8; // @[VCR.scala 191:22:@607.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waddr = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  wstate = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rstate = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  rdata = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_0 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_1 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_2 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_3 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_4 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_5 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_6 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_7 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  reg_8 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  reg_9 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      waddr <= 16'hffff;
    end else begin
      if (_T_162) begin
        waddr <= io_host_aw_bits_addr;
      end
    end
    if (reset) begin
      wstate <= 2'h0;
    end else begin
      if (_T_159) begin
        if (io_host_aw_valid) begin
          wstate <= 2'h1;
        end
      end else begin
        if (_T_160) begin
          if (io_host_w_valid) begin
            wstate <= 2'h2;
          end
        end else begin
          if (_T_161) begin
            if (io_host_b_ready) begin
              wstate <= 2'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      rstate <= 1'h0;
    end else begin
      if (_T_167) begin
        if (io_host_ar_valid) begin
          rstate <= 1'h1;
        end
      end else begin
        if (rstate) begin
          if (io_host_r_ready) begin
            rstate <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      rdata <= 32'h0;
    end else begin
      if (_T_209) begin
        if (_T_229) begin
          rdata <= reg_0;
        end else begin
          if (_T_227) begin
            rdata <= reg_1;
          end else begin
            if (_T_225) begin
              rdata <= reg_2;
            end else begin
              if (_T_223) begin
                rdata <= reg_3;
              end else begin
                if (_T_221) begin
                  rdata <= reg_4;
                end else begin
                  if (_T_219) begin
                    rdata <= reg_5;
                  end else begin
                    if (_T_217) begin
                      rdata <= reg_6;
                    end else begin
                      if (_T_215) begin
                        rdata <= reg_7;
                      end else begin
                        if (_T_213) begin
                          rdata <= reg_8;
                        end else begin
                          if (_T_211) begin
                            rdata <= reg_9;
                          end else begin
                            rdata <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_0 <= 32'h0;
    end else begin
      if (io_vcr_finish) begin
        reg_0 <= 32'h2;
      end else begin
        if (_T_176) begin
          reg_0 <= io_host_w_bits_data;
        end
      end
    end
    if (reset) begin
      reg_1 <= 32'h0;
    end else begin
      if (io_vcr_ecnt_0_valid) begin
        reg_1 <= io_vcr_ecnt_0_bits;
      end else begin
        if (_T_180) begin
          reg_1 <= io_host_w_bits_data;
        end
      end
    end
    if (reset) begin
      reg_2 <= 32'h0;
    end else begin
      if (_T_184) begin
        reg_2 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_3 <= 32'h0;
    end else begin
      if (_T_188) begin
        reg_3 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_4 <= 32'h0;
    end else begin
      if (_T_192) begin
        reg_4 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_5 <= 32'h0;
    end else begin
      if (_T_196) begin
        reg_5 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_6 <= 32'h0;
    end else begin
      if (_T_200) begin
        reg_6 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_7 <= 32'h0;
    end else begin
      if (_T_204) begin
        reg_7 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_8 <= 32'h0;
    end else begin
      if (_T_208) begin
        reg_8 <= io_host_w_bits_data;
      end
    end
    if (reset) begin
      reg_9 <= 32'h0;
    end else begin
      if (io_vcr_ucnt_0_valid) begin
        reg_9 <= io_vcr_ucnt_0_bits;
      end else begin
        if (_T_235) begin
          reg_9 <= io_host_w_bits_data;
        end
      end
    end
  end
endmodule
module Arbiter( // @[:@619.2]
  output        io_in_0_ready, // @[:@622.4]
  input         io_in_0_valid, // @[:@622.4]
  input  [31:0] io_in_0_bits_addr, // @[:@622.4]
  input  [7:0]  io_in_0_bits_len, // @[:@622.4]
  output        io_in_1_ready, // @[:@622.4]
  input         io_in_1_valid, // @[:@622.4]
  input  [31:0] io_in_1_bits_addr, // @[:@622.4]
  input  [7:0]  io_in_1_bits_len, // @[:@622.4]
  output        io_in_2_ready, // @[:@622.4]
  input         io_in_2_valid, // @[:@622.4]
  input  [31:0] io_in_2_bits_addr, // @[:@622.4]
  input  [7:0]  io_in_2_bits_len, // @[:@622.4]
  output        io_in_3_ready, // @[:@622.4]
  input         io_in_3_valid, // @[:@622.4]
  input  [31:0] io_in_3_bits_addr, // @[:@622.4]
  input  [7:0]  io_in_3_bits_len, // @[:@622.4]
  output        io_in_4_ready, // @[:@622.4]
  input         io_in_4_valid, // @[:@622.4]
  input  [31:0] io_in_4_bits_addr, // @[:@622.4]
  input  [7:0]  io_in_4_bits_len, // @[:@622.4]
  input         io_out_ready, // @[:@622.4]
  output        io_out_valid, // @[:@622.4]
  output [31:0] io_out_bits_addr, // @[:@622.4]
  output [7:0]  io_out_bits_len, // @[:@622.4]
  output [2:0]  io_chosen // @[:@622.4]
);
  wire [2:0] _GEN_0; // @[Arbiter.scala 126:27:@627.4]
  wire [7:0] _GEN_1; // @[Arbiter.scala 126:27:@627.4]
  wire [31:0] _GEN_2; // @[Arbiter.scala 126:27:@627.4]
  wire [2:0] _GEN_3; // @[Arbiter.scala 126:27:@632.4]
  wire [7:0] _GEN_4; // @[Arbiter.scala 126:27:@632.4]
  wire [31:0] _GEN_5; // @[Arbiter.scala 126:27:@632.4]
  wire [2:0] _GEN_6; // @[Arbiter.scala 126:27:@637.4]
  wire [7:0] _GEN_7; // @[Arbiter.scala 126:27:@637.4]
  wire [31:0] _GEN_8; // @[Arbiter.scala 126:27:@637.4]
  wire  _T_114; // @[Arbiter.scala 31:68:@647.4]
  wire  _T_115; // @[Arbiter.scala 31:68:@648.4]
  wire  _T_116; // @[Arbiter.scala 31:68:@649.4]
  wire  _T_118; // @[Arbiter.scala 31:78:@650.4]
  wire  _T_120; // @[Arbiter.scala 31:78:@651.4]
  wire  _T_122; // @[Arbiter.scala 31:78:@652.4]
  wire  _T_124; // @[Arbiter.scala 31:78:@653.4]
  wire  _T_131; // @[Arbiter.scala 135:19:@664.4]
  assign _GEN_0 = io_in_3_valid ? 3'h3 : 3'h4; // @[Arbiter.scala 126:27:@627.4]
  assign _GEN_1 = io_in_3_valid ? io_in_3_bits_len : io_in_4_bits_len; // @[Arbiter.scala 126:27:@627.4]
  assign _GEN_2 = io_in_3_valid ? io_in_3_bits_addr : io_in_4_bits_addr; // @[Arbiter.scala 126:27:@627.4]
  assign _GEN_3 = io_in_2_valid ? 3'h2 : _GEN_0; // @[Arbiter.scala 126:27:@632.4]
  assign _GEN_4 = io_in_2_valid ? io_in_2_bits_len : _GEN_1; // @[Arbiter.scala 126:27:@632.4]
  assign _GEN_5 = io_in_2_valid ? io_in_2_bits_addr : _GEN_2; // @[Arbiter.scala 126:27:@632.4]
  assign _GEN_6 = io_in_1_valid ? 3'h1 : _GEN_3; // @[Arbiter.scala 126:27:@637.4]
  assign _GEN_7 = io_in_1_valid ? io_in_1_bits_len : _GEN_4; // @[Arbiter.scala 126:27:@637.4]
  assign _GEN_8 = io_in_1_valid ? io_in_1_bits_addr : _GEN_5; // @[Arbiter.scala 126:27:@637.4]
  assign _T_114 = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68:@647.4]
  assign _T_115 = _T_114 | io_in_2_valid; // @[Arbiter.scala 31:68:@648.4]
  assign _T_116 = _T_115 | io_in_3_valid; // @[Arbiter.scala 31:68:@649.4]
  assign _T_118 = io_in_0_valid == 1'h0; // @[Arbiter.scala 31:78:@650.4]
  assign _T_120 = _T_114 == 1'h0; // @[Arbiter.scala 31:78:@651.4]
  assign _T_122 = _T_115 == 1'h0; // @[Arbiter.scala 31:78:@652.4]
  assign _T_124 = _T_116 == 1'h0; // @[Arbiter.scala 31:78:@653.4]
  assign _T_131 = _T_124 == 1'h0; // @[Arbiter.scala 135:19:@664.4]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14:@655.4]
  assign io_in_1_ready = _T_118 & io_out_ready; // @[Arbiter.scala 134:14:@657.4]
  assign io_in_2_ready = _T_120 & io_out_ready; // @[Arbiter.scala 134:14:@659.4]
  assign io_in_3_ready = _T_122 & io_out_ready; // @[Arbiter.scala 134:14:@661.4]
  assign io_in_4_ready = _T_124 & io_out_ready; // @[Arbiter.scala 134:14:@663.4]
  assign io_out_valid = _T_131 | io_in_4_valid; // @[Arbiter.scala 135:16:@666.4]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_8; // @[Arbiter.scala 124:15:@626.4 Arbiter.scala 128:19:@630.6 Arbiter.scala 128:19:@635.6 Arbiter.scala 128:19:@640.6 Arbiter.scala 128:19:@645.6]
  assign io_out_bits_len = io_in_0_valid ? io_in_0_bits_len : _GEN_7; // @[Arbiter.scala 124:15:@625.4 Arbiter.scala 128:19:@629.6 Arbiter.scala 128:19:@634.6 Arbiter.scala 128:19:@639.6 Arbiter.scala 128:19:@644.6]
  assign io_chosen = io_in_0_valid ? 3'h0 : _GEN_6; // @[Arbiter.scala 123:13:@624.4 Arbiter.scala 127:17:@628.6 Arbiter.scala 127:17:@633.6 Arbiter.scala 127:17:@638.6 Arbiter.scala 127:17:@643.6]
endmodule
module VME( // @[:@668.2]
  input         clock, // @[:@669.4]
  input         reset, // @[:@670.4]
  input         io_mem_aw_ready, // @[:@671.4]
  output        io_mem_aw_valid, // @[:@671.4]
  output [31:0] io_mem_aw_bits_addr, // @[:@671.4]
  output [7:0]  io_mem_aw_bits_len, // @[:@671.4]
  input         io_mem_w_ready, // @[:@671.4]
  output        io_mem_w_valid, // @[:@671.4]
  output [63:0] io_mem_w_bits_data, // @[:@671.4]
  output        io_mem_w_bits_last, // @[:@671.4]
  output        io_mem_b_ready, // @[:@671.4]
  input         io_mem_b_valid, // @[:@671.4]
  input         io_mem_ar_ready, // @[:@671.4]
  output        io_mem_ar_valid, // @[:@671.4]
  output [31:0] io_mem_ar_bits_addr, // @[:@671.4]
  output [7:0]  io_mem_ar_bits_len, // @[:@671.4]
  output        io_mem_r_ready, // @[:@671.4]
  input         io_mem_r_valid, // @[:@671.4]
  input  [63:0] io_mem_r_bits_data, // @[:@671.4]
  input         io_mem_r_bits_last, // @[:@671.4]
  output        io_vme_rd_0_cmd_ready, // @[:@671.4]
  input         io_vme_rd_0_cmd_valid, // @[:@671.4]
  input  [31:0] io_vme_rd_0_cmd_bits_addr, // @[:@671.4]
  input  [7:0]  io_vme_rd_0_cmd_bits_len, // @[:@671.4]
  input         io_vme_rd_0_data_ready, // @[:@671.4]
  output        io_vme_rd_0_data_valid, // @[:@671.4]
  output [63:0] io_vme_rd_0_data_bits, // @[:@671.4]
  output        io_vme_rd_1_cmd_ready, // @[:@671.4]
  input         io_vme_rd_1_cmd_valid, // @[:@671.4]
  input  [31:0] io_vme_rd_1_cmd_bits_addr, // @[:@671.4]
  input  [7:0]  io_vme_rd_1_cmd_bits_len, // @[:@671.4]
  input         io_vme_rd_1_data_ready, // @[:@671.4]
  output        io_vme_rd_1_data_valid, // @[:@671.4]
  output [63:0] io_vme_rd_1_data_bits, // @[:@671.4]
  output        io_vme_rd_2_cmd_ready, // @[:@671.4]
  input         io_vme_rd_2_cmd_valid, // @[:@671.4]
  input  [31:0] io_vme_rd_2_cmd_bits_addr, // @[:@671.4]
  input  [7:0]  io_vme_rd_2_cmd_bits_len, // @[:@671.4]
  input         io_vme_rd_2_data_ready, // @[:@671.4]
  output        io_vme_rd_2_data_valid, // @[:@671.4]
  output [63:0] io_vme_rd_2_data_bits, // @[:@671.4]
  output        io_vme_rd_3_cmd_ready, // @[:@671.4]
  input         io_vme_rd_3_cmd_valid, // @[:@671.4]
  input  [31:0] io_vme_rd_3_cmd_bits_addr, // @[:@671.4]
  input  [7:0]  io_vme_rd_3_cmd_bits_len, // @[:@671.4]
  input         io_vme_rd_3_data_ready, // @[:@671.4]
  output        io_vme_rd_3_data_valid, // @[:@671.4]
  output [63:0] io_vme_rd_3_data_bits, // @[:@671.4]
  output        io_vme_rd_4_cmd_ready, // @[:@671.4]
  input         io_vme_rd_4_cmd_valid, // @[:@671.4]
  input  [31:0] io_vme_rd_4_cmd_bits_addr, // @[:@671.4]
  input  [7:0]  io_vme_rd_4_cmd_bits_len, // @[:@671.4]
  input         io_vme_rd_4_data_ready, // @[:@671.4]
  output        io_vme_rd_4_data_valid, // @[:@671.4]
  output [63:0] io_vme_rd_4_data_bits, // @[:@671.4]
  output        io_vme_wr_0_cmd_ready, // @[:@671.4]
  input         io_vme_wr_0_cmd_valid, // @[:@671.4]
  input  [31:0] io_vme_wr_0_cmd_bits_addr, // @[:@671.4]
  input  [7:0]  io_vme_wr_0_cmd_bits_len, // @[:@671.4]
  output        io_vme_wr_0_data_ready, // @[:@671.4]
  input         io_vme_wr_0_data_valid, // @[:@671.4]
  input  [63:0] io_vme_wr_0_data_bits, // @[:@671.4]
  output        io_vme_wr_0_ack // @[:@671.4]
);
  wire  rd_arb_io_in_0_ready; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_in_0_valid; // @[VME.scala 146:22:@673.4]
  wire [31:0] rd_arb_io_in_0_bits_addr; // @[VME.scala 146:22:@673.4]
  wire [7:0] rd_arb_io_in_0_bits_len; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_in_1_ready; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_in_1_valid; // @[VME.scala 146:22:@673.4]
  wire [31:0] rd_arb_io_in_1_bits_addr; // @[VME.scala 146:22:@673.4]
  wire [7:0] rd_arb_io_in_1_bits_len; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_in_2_ready; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_in_2_valid; // @[VME.scala 146:22:@673.4]
  wire [31:0] rd_arb_io_in_2_bits_addr; // @[VME.scala 146:22:@673.4]
  wire [7:0] rd_arb_io_in_2_bits_len; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_in_3_ready; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_in_3_valid; // @[VME.scala 146:22:@673.4]
  wire [31:0] rd_arb_io_in_3_bits_addr; // @[VME.scala 146:22:@673.4]
  wire [7:0] rd_arb_io_in_3_bits_len; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_in_4_ready; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_in_4_valid; // @[VME.scala 146:22:@673.4]
  wire [31:0] rd_arb_io_in_4_bits_addr; // @[VME.scala 146:22:@673.4]
  wire [7:0] rd_arb_io_in_4_bits_len; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_out_ready; // @[VME.scala 146:22:@673.4]
  wire  rd_arb_io_out_valid; // @[VME.scala 146:22:@673.4]
  wire [31:0] rd_arb_io_out_bits_addr; // @[VME.scala 146:22:@673.4]
  wire [7:0] rd_arb_io_out_bits_len; // @[VME.scala 146:22:@673.4]
  wire [2:0] rd_arb_io_chosen; // @[VME.scala 146:22:@673.4]
  wire  _T_260; // @[Decoupled.scala 37:37:@676.4]
  reg [2:0] rd_arb_chosen; // @[Reg.scala 11:16:@677.4]
  reg [31:0] _RAND_0;
  reg [1:0] rstate; // @[VME.scala 152:23:@701.4]
  reg [31:0] _RAND_1;
  wire  _T_263; // @[Conditional.scala 37:30:@702.4]
  wire [1:0] _GEN_1; // @[VME.scala 156:33:@704.6]
  wire  _T_264; // @[Conditional.scala 37:30:@709.6]
  wire [1:0] _GEN_2; // @[VME.scala 161:29:@711.8]
  wire  _T_265; // @[Conditional.scala 37:30:@716.8]
  wire  _T_266; // @[Decoupled.scala 37:37:@718.10]
  wire  _T_267; // @[VME.scala 166:28:@719.10]
  wire [1:0] _GEN_3; // @[VME.scala 166:51:@720.10]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@717.8]
  wire [1:0] _GEN_5; // @[Conditional.scala 39:67:@710.6]
  wire [1:0] _GEN_6; // @[Conditional.scala 40:58:@703.4]
  reg [1:0] wstate; // @[VME.scala 173:23:@724.4]
  reg [31:0] _RAND_2;
  reg [7:0] wr_cnt; // @[VME.scala 176:23:@725.4]
  reg [31:0] _RAND_3;
  wire  _T_271; // @[VME.scala 178:15:@726.4]
  wire  _T_273; // @[Decoupled.scala 37:37:@731.6]
  wire [8:0] _T_275; // @[VME.scala 181:22:@733.8]
  wire [7:0] _T_276; // @[VME.scala 181:22:@734.8]
  wire [7:0] _GEN_7; // @[VME.scala 180:31:@732.6]
  wire [7:0] _GEN_8; // @[VME.scala 178:31:@727.4]
  wire  _T_277; // @[Conditional.scala 37:30:@737.4]
  wire [1:0] _GEN_9; // @[VME.scala 186:36:@739.6]
  wire  _T_278; // @[Conditional.scala 37:30:@744.6]
  wire [1:0] _GEN_10; // @[VME.scala 191:29:@746.8]
  wire  _T_279; // @[Conditional.scala 37:30:@751.8]
  wire  _T_280; // @[VME.scala 200:18:@753.10]
  wire  _T_281; // @[VME.scala 200:46:@754.10]
  wire  _T_282; // @[VME.scala 200:36:@755.10]
  wire [1:0] _GEN_11; // @[VME.scala 200:77:@756.10]
  wire  _T_283; // @[Conditional.scala 37:30:@761.10]
  wire [1:0] _GEN_12; // @[VME.scala 205:28:@763.12]
  wire [1:0] _GEN_13; // @[Conditional.scala 39:67:@762.10]
  wire [1:0] _GEN_14; // @[Conditional.scala 39:67:@752.8]
  wire [1:0] _GEN_15; // @[Conditional.scala 39:67:@745.6]
  wire [1:0] _GEN_16; // @[Conditional.scala 40:58:@738.4]
  reg [7:0] rd_len; // @[VME.scala 213:23:@767.4]
  reg [31:0] _RAND_4;
  reg [7:0] wr_len; // @[VME.scala 214:23:@768.4]
  reg [31:0] _RAND_5;
  reg [31:0] rd_addr; // @[VME.scala 215:24:@769.4]
  reg [31:0] _RAND_6;
  reg [31:0] wr_addr; // @[VME.scala 216:24:@770.4]
  reg [31:0] _RAND_7;
  wire [7:0] _GEN_17; // @[VME.scala 218:30:@772.4]
  wire [31:0] _GEN_18; // @[VME.scala 218:30:@772.4]
  wire  _T_293; // @[Decoupled.scala 37:37:@776.4]
  wire [7:0] _GEN_19; // @[VME.scala 223:33:@777.4]
  wire [31:0] _GEN_20; // @[VME.scala 223:33:@777.4]
  wire  _T_296; // @[VME.scala 233:46:@783.4]
  wire  _T_299; // @[VME.scala 233:46:@787.4]
  wire  _T_302; // @[VME.scala 233:46:@791.4]
  wire  _T_305; // @[VME.scala 233:46:@795.4]
  wire  _T_308; // @[VME.scala 233:46:@799.4]
  wire  _T_312; // @[VME.scala 239:37:@807.4]
  wire  _T_320; // @[VME.scala 256:28:@826.4]
  wire  _GEN_32; // @[VME.scala 256:42:@827.4]
  wire  _GEN_39; // @[VME.scala 256:42:@827.4]
  wire  _GEN_46; // @[VME.scala 256:42:@827.4]
  wire  _GEN_53; // @[VME.scala 256:42:@827.4]
  Arbiter rd_arb ( // @[VME.scala 146:22:@673.4]
    .io_in_0_ready(rd_arb_io_in_0_ready),
    .io_in_0_valid(rd_arb_io_in_0_valid),
    .io_in_0_bits_addr(rd_arb_io_in_0_bits_addr),
    .io_in_0_bits_len(rd_arb_io_in_0_bits_len),
    .io_in_1_ready(rd_arb_io_in_1_ready),
    .io_in_1_valid(rd_arb_io_in_1_valid),
    .io_in_1_bits_addr(rd_arb_io_in_1_bits_addr),
    .io_in_1_bits_len(rd_arb_io_in_1_bits_len),
    .io_in_2_ready(rd_arb_io_in_2_ready),
    .io_in_2_valid(rd_arb_io_in_2_valid),
    .io_in_2_bits_addr(rd_arb_io_in_2_bits_addr),
    .io_in_2_bits_len(rd_arb_io_in_2_bits_len),
    .io_in_3_ready(rd_arb_io_in_3_ready),
    .io_in_3_valid(rd_arb_io_in_3_valid),
    .io_in_3_bits_addr(rd_arb_io_in_3_bits_addr),
    .io_in_3_bits_len(rd_arb_io_in_3_bits_len),
    .io_in_4_ready(rd_arb_io_in_4_ready),
    .io_in_4_valid(rd_arb_io_in_4_valid),
    .io_in_4_bits_addr(rd_arb_io_in_4_bits_addr),
    .io_in_4_bits_len(rd_arb_io_in_4_bits_len),
    .io_out_ready(rd_arb_io_out_ready),
    .io_out_valid(rd_arb_io_out_valid),
    .io_out_bits_addr(rd_arb_io_out_bits_addr),
    .io_out_bits_len(rd_arb_io_out_bits_len),
    .io_chosen(rd_arb_io_chosen)
  );
  assign _T_260 = rd_arb_io_out_ready & rd_arb_io_out_valid; // @[Decoupled.scala 37:37:@676.4]
  assign _T_263 = 2'h0 == rstate; // @[Conditional.scala 37:30:@702.4]
  assign _GEN_1 = rd_arb_io_out_valid ? 2'h1 : rstate; // @[VME.scala 156:33:@704.6]
  assign _T_264 = 2'h1 == rstate; // @[Conditional.scala 37:30:@709.6]
  assign _GEN_2 = io_mem_ar_ready ? 2'h2 : rstate; // @[VME.scala 161:29:@711.8]
  assign _T_265 = 2'h2 == rstate; // @[Conditional.scala 37:30:@716.8]
  assign _T_266 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 37:37:@718.10]
  assign _T_267 = _T_266 & io_mem_r_bits_last; // @[VME.scala 166:28:@719.10]
  assign _GEN_3 = _T_267 ? 2'h0 : rstate; // @[VME.scala 166:51:@720.10]
  assign _GEN_4 = _T_265 ? _GEN_3 : rstate; // @[Conditional.scala 39:67:@717.8]
  assign _GEN_5 = _T_264 ? _GEN_2 : _GEN_4; // @[Conditional.scala 39:67:@710.6]
  assign _GEN_6 = _T_263 ? _GEN_1 : _GEN_5; // @[Conditional.scala 40:58:@703.4]
  assign _T_271 = wstate == 2'h0; // @[VME.scala 178:15:@726.4]
  assign _T_273 = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 37:37:@731.6]
  assign _T_275 = wr_cnt + 8'h1; // @[VME.scala 181:22:@733.8]
  assign _T_276 = wr_cnt + 8'h1; // @[VME.scala 181:22:@734.8]
  assign _GEN_7 = _T_273 ? _T_276 : wr_cnt; // @[VME.scala 180:31:@732.6]
  assign _GEN_8 = _T_271 ? 8'h0 : _GEN_7; // @[VME.scala 178:31:@727.4]
  assign _T_277 = 2'h0 == wstate; // @[Conditional.scala 37:30:@737.4]
  assign _GEN_9 = io_vme_wr_0_cmd_valid ? 2'h1 : wstate; // @[VME.scala 186:36:@739.6]
  assign _T_278 = 2'h1 == wstate; // @[Conditional.scala 37:30:@744.6]
  assign _GEN_10 = io_mem_aw_ready ? 2'h2 : wstate; // @[VME.scala 191:29:@746.8]
  assign _T_279 = 2'h2 == wstate; // @[Conditional.scala 37:30:@751.8]
  assign _T_280 = io_vme_wr_0_data_valid & io_mem_w_ready; // @[VME.scala 200:18:@753.10]
  assign _T_281 = wr_cnt == io_vme_wr_0_cmd_bits_len; // @[VME.scala 200:46:@754.10]
  assign _T_282 = _T_280 & _T_281; // @[VME.scala 200:36:@755.10]
  assign _GEN_11 = _T_282 ? 2'h3 : wstate; // @[VME.scala 200:77:@756.10]
  assign _T_283 = 2'h3 == wstate; // @[Conditional.scala 37:30:@761.10]
  assign _GEN_12 = io_mem_b_valid ? 2'h0 : wstate; // @[VME.scala 205:28:@763.12]
  assign _GEN_13 = _T_283 ? _GEN_12 : wstate; // @[Conditional.scala 39:67:@762.10]
  assign _GEN_14 = _T_279 ? _GEN_11 : _GEN_13; // @[Conditional.scala 39:67:@752.8]
  assign _GEN_15 = _T_278 ? _GEN_10 : _GEN_14; // @[Conditional.scala 39:67:@745.6]
  assign _GEN_16 = _T_277 ? _GEN_9 : _GEN_15; // @[Conditional.scala 40:58:@738.4]
  assign _GEN_17 = _T_260 ? rd_arb_io_out_bits_len : rd_len; // @[VME.scala 218:30:@772.4]
  assign _GEN_18 = _T_260 ? rd_arb_io_out_bits_addr : rd_addr; // @[VME.scala 218:30:@772.4]
  assign _T_293 = io_vme_wr_0_cmd_ready & io_vme_wr_0_cmd_valid; // @[Decoupled.scala 37:37:@776.4]
  assign _GEN_19 = _T_293 ? io_vme_wr_0_cmd_bits_len : wr_len; // @[VME.scala 223:33:@777.4]
  assign _GEN_20 = _T_293 ? io_vme_wr_0_cmd_bits_addr : wr_addr; // @[VME.scala 223:33:@777.4]
  assign _T_296 = rd_arb_chosen == 3'h0; // @[VME.scala 233:46:@783.4]
  assign _T_299 = rd_arb_chosen == 3'h1; // @[VME.scala 233:46:@787.4]
  assign _T_302 = rd_arb_chosen == 3'h2; // @[VME.scala 233:46:@791.4]
  assign _T_305 = rd_arb_chosen == 3'h3; // @[VME.scala 233:46:@795.4]
  assign _T_308 = rd_arb_chosen == 3'h4; // @[VME.scala 233:46:@799.4]
  assign _T_312 = wstate == 2'h2; // @[VME.scala 239:37:@807.4]
  assign _T_320 = rstate == 2'h2; // @[VME.scala 256:28:@826.4]
  assign _GEN_32 = 3'h1 == rd_arb_chosen ? io_vme_rd_1_data_ready : io_vme_rd_0_data_ready; // @[VME.scala 256:42:@827.4]
  assign _GEN_39 = 3'h2 == rd_arb_chosen ? io_vme_rd_2_data_ready : _GEN_32; // @[VME.scala 256:42:@827.4]
  assign _GEN_46 = 3'h3 == rd_arb_chosen ? io_vme_rd_3_data_ready : _GEN_39; // @[VME.scala 256:42:@827.4]
  assign _GEN_53 = 3'h4 == rd_arb_chosen ? io_vme_rd_4_data_ready : _GEN_46; // @[VME.scala 256:42:@827.4]
  assign io_mem_aw_valid = wstate == 2'h1; // @[VME.scala 242:19:@811.4]
  assign io_mem_aw_bits_addr = wr_addr; // @[VME.scala 243:23:@812.4]
  assign io_mem_aw_bits_len = wr_len; // @[VME.scala 244:22:@813.4]
  assign io_mem_w_valid = _T_312 & io_vme_wr_0_data_valid; // @[VME.scala 246:18:@816.4]
  assign io_mem_w_bits_data = io_vme_wr_0_data_bits; // @[VME.scala 247:22:@817.4]
  assign io_mem_w_bits_last = wr_cnt == io_vme_wr_0_cmd_bits_len; // @[VME.scala 248:22:@819.4]
  assign io_mem_b_ready = wstate == 2'h3; // @[VME.scala 250:18:@821.4]
  assign io_mem_ar_valid = rstate == 2'h1; // @[VME.scala 252:19:@823.4]
  assign io_mem_ar_bits_addr = rd_addr; // @[VME.scala 253:23:@824.4]
  assign io_mem_ar_bits_len = rd_len; // @[VME.scala 254:22:@825.4]
  assign io_mem_r_ready = _T_320 & _GEN_53; // @[VME.scala 256:18:@828.4]
  assign io_vme_rd_0_cmd_ready = rd_arb_io_in_0_ready; // @[VME.scala 149:53:@684.4]
  assign io_vme_rd_0_data_valid = _T_296 & io_mem_r_valid; // @[VME.scala 233:29:@785.4]
  assign io_vme_rd_0_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@786.4]
  assign io_vme_rd_1_cmd_ready = rd_arb_io_in_1_ready; // @[VME.scala 149:53:@688.4]
  assign io_vme_rd_1_data_valid = _T_299 & io_mem_r_valid; // @[VME.scala 233:29:@789.4]
  assign io_vme_rd_1_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@790.4]
  assign io_vme_rd_2_cmd_ready = rd_arb_io_in_2_ready; // @[VME.scala 149:53:@692.4]
  assign io_vme_rd_2_data_valid = _T_302 & io_mem_r_valid; // @[VME.scala 233:29:@793.4]
  assign io_vme_rd_2_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@794.4]
  assign io_vme_rd_3_cmd_ready = rd_arb_io_in_3_ready; // @[VME.scala 149:53:@696.4]
  assign io_vme_rd_3_data_valid = _T_305 & io_mem_r_valid; // @[VME.scala 233:29:@797.4]
  assign io_vme_rd_3_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@798.4]
  assign io_vme_rd_4_cmd_ready = rd_arb_io_in_4_ready; // @[VME.scala 149:53:@700.4]
  assign io_vme_rd_4_data_valid = _T_308 & io_mem_r_valid; // @[VME.scala 233:29:@801.4]
  assign io_vme_rd_4_data_bits = io_mem_r_bits_data; // @[VME.scala 234:28:@802.4]
  assign io_vme_wr_0_cmd_ready = wstate == 2'h0; // @[VME.scala 237:26:@804.4]
  assign io_vme_wr_0_data_ready = _T_312 & io_mem_w_ready; // @[VME.scala 239:27:@809.4]
  assign io_vme_wr_0_ack = io_mem_b_ready & io_mem_b_valid; // @[VME.scala 238:20:@806.4]
  assign rd_arb_io_in_0_valid = io_vme_rd_0_cmd_valid; // @[VME.scala 149:53:@683.4]
  assign rd_arb_io_in_0_bits_addr = io_vme_rd_0_cmd_bits_addr; // @[VME.scala 149:53:@682.4]
  assign rd_arb_io_in_0_bits_len = io_vme_rd_0_cmd_bits_len; // @[VME.scala 149:53:@681.4]
  assign rd_arb_io_in_1_valid = io_vme_rd_1_cmd_valid; // @[VME.scala 149:53:@687.4]
  assign rd_arb_io_in_1_bits_addr = io_vme_rd_1_cmd_bits_addr; // @[VME.scala 149:53:@686.4]
  assign rd_arb_io_in_1_bits_len = io_vme_rd_1_cmd_bits_len; // @[VME.scala 149:53:@685.4]
  assign rd_arb_io_in_2_valid = io_vme_rd_2_cmd_valid; // @[VME.scala 149:53:@691.4]
  assign rd_arb_io_in_2_bits_addr = io_vme_rd_2_cmd_bits_addr; // @[VME.scala 149:53:@690.4]
  assign rd_arb_io_in_2_bits_len = io_vme_rd_2_cmd_bits_len; // @[VME.scala 149:53:@689.4]
  assign rd_arb_io_in_3_valid = io_vme_rd_3_cmd_valid; // @[VME.scala 149:53:@695.4]
  assign rd_arb_io_in_3_bits_addr = io_vme_rd_3_cmd_bits_addr; // @[VME.scala 149:53:@694.4]
  assign rd_arb_io_in_3_bits_len = io_vme_rd_3_cmd_bits_len; // @[VME.scala 149:53:@693.4]
  assign rd_arb_io_in_4_valid = io_vme_rd_4_cmd_valid; // @[VME.scala 149:53:@699.4]
  assign rd_arb_io_in_4_bits_addr = io_vme_rd_4_cmd_bits_addr; // @[VME.scala 149:53:@698.4]
  assign rd_arb_io_in_4_bits_len = io_vme_rd_4_cmd_bits_len; // @[VME.scala 149:53:@697.4]
  assign rd_arb_io_out_ready = rstate == 2'h0; // @[VME.scala 229:23:@782.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_arb_chosen = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rstate = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  wstate = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  wr_cnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_len = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  wr_len = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  wr_addr = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_260) begin
      rd_arb_chosen <= rd_arb_io_chosen;
    end
    if (reset) begin
      rstate <= 2'h0;
    end else begin
      if (_T_263) begin
        if (rd_arb_io_out_valid) begin
          rstate <= 2'h1;
        end
      end else begin
        if (_T_264) begin
          if (io_mem_ar_ready) begin
            rstate <= 2'h2;
          end
        end else begin
          if (_T_265) begin
            if (_T_267) begin
              rstate <= 2'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      wstate <= 2'h0;
    end else begin
      if (_T_277) begin
        if (io_vme_wr_0_cmd_valid) begin
          wstate <= 2'h1;
        end
      end else begin
        if (_T_278) begin
          if (io_mem_aw_ready) begin
            wstate <= 2'h2;
          end
        end else begin
          if (_T_279) begin
            if (_T_282) begin
              wstate <= 2'h3;
            end
          end else begin
            if (_T_283) begin
              if (io_mem_b_valid) begin
                wstate <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      wr_cnt <= 8'h0;
    end else begin
      if (_T_271) begin
        wr_cnt <= 8'h0;
      end else begin
        if (_T_273) begin
          wr_cnt <= _T_276;
        end
      end
    end
    if (reset) begin
      rd_len <= 8'h0;
    end else begin
      if (_T_260) begin
        rd_len <= rd_arb_io_out_bits_len;
      end
    end
    if (reset) begin
      wr_len <= 8'h0;
    end else begin
      if (_T_293) begin
        wr_len <= io_vme_wr_0_cmd_bits_len;
      end
    end
    if (reset) begin
      rd_addr <= 32'h0;
    end else begin
      if (_T_260) begin
        rd_addr <= rd_arb_io_out_bits_addr;
      end
    end
    if (reset) begin
      wr_addr <= 32'h0;
    end else begin
      if (_T_293) begin
        wr_addr <= io_vme_wr_0_cmd_bits_addr;
      end
    end
  end
endmodule
module Queue( // @[:@852.2]
  input          clock, // @[:@853.4]
  input          reset, // @[:@854.4]
  output         io_enq_ready, // @[:@855.4]
  input          io_enq_valid, // @[:@855.4]
  input  [127:0] io_enq_bits, // @[:@855.4]
  input          io_deq_ready, // @[:@855.4]
  output         io_deq_valid, // @[:@855.4]
  output [127:0] io_deq_bits, // @[:@855.4]
  output [7:0]   io_count // @[:@855.4]
);
  reg [127:0] _T_35 [0:127]; // @[Decoupled.scala 215:24:@857.4]
  reg [127:0] _RAND_0;
  wire [127:0] _T_35__T_68_data; // @[Decoupled.scala 215:24:@857.4]
  wire [6:0] _T_35__T_68_addr; // @[Decoupled.scala 215:24:@857.4]
  wire [127:0] _T_35__T_54_data; // @[Decoupled.scala 215:24:@857.4]
  wire [6:0] _T_35__T_54_addr; // @[Decoupled.scala 215:24:@857.4]
  wire  _T_35__T_54_mask; // @[Decoupled.scala 215:24:@857.4]
  wire  _T_35__T_54_en; // @[Decoupled.scala 215:24:@857.4]
  reg [6:0] value; // @[Counter.scala 26:33:@858.4]
  reg [31:0] _RAND_1;
  reg [6:0] value_1; // @[Counter.scala 26:33:@859.4]
  reg [31:0] _RAND_2;
  reg  _T_42; // @[Decoupled.scala 218:35:@860.4]
  reg [31:0] _RAND_3;
  wire  _T_43; // @[Decoupled.scala 220:41:@861.4]
  wire  _T_45; // @[Decoupled.scala 221:36:@862.4]
  wire  _T_46; // @[Decoupled.scala 221:33:@863.4]
  wire  _T_47; // @[Decoupled.scala 222:32:@864.4]
  wire  _T_48; // @[Decoupled.scala 37:37:@865.4]
  wire  _T_51; // @[Decoupled.scala 37:37:@868.4]
  wire [7:0] _T_57; // @[Counter.scala 35:22:@875.6]
  wire [6:0] _T_58; // @[Counter.scala 35:22:@876.6]
  wire [6:0] _GEN_5; // @[Decoupled.scala 226:17:@871.4]
  wire [7:0] _T_61; // @[Counter.scala 35:22:@881.6]
  wire [6:0] _T_62; // @[Counter.scala 35:22:@882.6]
  wire [6:0] _GEN_6; // @[Decoupled.scala 230:17:@879.4]
  wire  _T_63; // @[Decoupled.scala 233:16:@885.4]
  wire  _GEN_7; // @[Decoupled.scala 233:28:@886.4]
  wire [7:0] _T_69; // @[Decoupled.scala 254:40:@895.4]
  wire [7:0] _T_70; // @[Decoupled.scala 254:40:@896.4]
  wire [6:0] _T_71; // @[Decoupled.scala 254:40:@897.4]
  wire  _T_72; // @[Decoupled.scala 256:32:@898.4]
  wire [7:0] _T_75; // @[Decoupled.scala 256:20:@899.4]
  wire [7:0] _GEN_14; // @[Decoupled.scala 256:62:@900.4]
  assign _T_35__T_68_addr = value_1;
  assign _T_35__T_68_data = _T_35[_T_35__T_68_addr]; // @[Decoupled.scala 215:24:@857.4]
  assign _T_35__T_54_data = io_enq_bits;
  assign _T_35__T_54_addr = value;
  assign _T_35__T_54_mask = 1'h1;
  assign _T_35__T_54_en = io_enq_ready & io_enq_valid;
  assign _T_43 = value == value_1; // @[Decoupled.scala 220:41:@861.4]
  assign _T_45 = _T_42 == 1'h0; // @[Decoupled.scala 221:36:@862.4]
  assign _T_46 = _T_43 & _T_45; // @[Decoupled.scala 221:33:@863.4]
  assign _T_47 = _T_43 & _T_42; // @[Decoupled.scala 222:32:@864.4]
  assign _T_48 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:@865.4]
  assign _T_51 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:@868.4]
  assign _T_57 = value + 7'h1; // @[Counter.scala 35:22:@875.6]
  assign _T_58 = value + 7'h1; // @[Counter.scala 35:22:@876.6]
  assign _GEN_5 = _T_48 ? _T_58 : value; // @[Decoupled.scala 226:17:@871.4]
  assign _T_61 = value_1 + 7'h1; // @[Counter.scala 35:22:@881.6]
  assign _T_62 = value_1 + 7'h1; // @[Counter.scala 35:22:@882.6]
  assign _GEN_6 = _T_51 ? _T_62 : value_1; // @[Decoupled.scala 230:17:@879.4]
  assign _T_63 = _T_48 != _T_51; // @[Decoupled.scala 233:16:@885.4]
  assign _GEN_7 = _T_63 ? _T_48 : _T_42; // @[Decoupled.scala 233:28:@886.4]
  assign _T_69 = value - value_1; // @[Decoupled.scala 254:40:@895.4]
  assign _T_70 = $unsigned(_T_69); // @[Decoupled.scala 254:40:@896.4]
  assign _T_71 = _T_70[6:0]; // @[Decoupled.scala 254:40:@897.4]
  assign _T_72 = _T_42 & _T_43; // @[Decoupled.scala 256:32:@898.4]
  assign _T_75 = _T_72 ? 8'h80 : 8'h0; // @[Decoupled.scala 256:20:@899.4]
  assign _GEN_14 = {{1'd0}, _T_71}; // @[Decoupled.scala 256:62:@900.4]
  assign io_enq_ready = _T_47 == 1'h0; // @[Decoupled.scala 238:16:@892.4]
  assign io_deq_valid = _T_46 == 1'h0; // @[Decoupled.scala 237:16:@890.4]
  assign io_deq_bits = _T_35__T_68_data; // @[Decoupled.scala 239:15:@894.4]
  assign io_count = _T_75 | _GEN_14; // @[Decoupled.scala 256:14:@901.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T_35[initvar] = _RAND_0[127:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_42 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35__T_54_en & _T_35__T_54_mask) begin
      _T_35[_T_35__T_54_addr] <= _T_35__T_54_data; // @[Decoupled.scala 215:24:@857.4]
    end
    if (reset) begin
      value <= 7'h0;
    end else begin
      if (_T_48) begin
        value <= _T_58;
      end
    end
    if (reset) begin
      value_1 <= 7'h0;
    end else begin
      if (_T_51) begin
        value_1 <= _T_62;
      end
    end
    if (reset) begin
      _T_42 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_42 <= _T_48;
      end
    end
  end
endmodule
module FetchDecode( // @[:@903.2]
  input  [127:0] io_inst, // @[:@906.4]
  output         io_isLoad, // @[:@906.4]
  output         io_isCompute, // @[:@906.4]
  output         io_isStore // @[:@906.4]
);
  wire [127:0] _T_15; // @[Lookup.scala 9:38:@908.4]
  wire  _T_16; // @[Lookup.scala 9:38:@909.4]
  wire  _T_20; // @[Lookup.scala 9:38:@911.4]
  wire  _T_24; // @[Lookup.scala 9:38:@913.4]
  wire  _T_28; // @[Lookup.scala 9:38:@915.4]
  wire [127:0] _T_31; // @[Lookup.scala 9:38:@916.4]
  wire  _T_32; // @[Lookup.scala 9:38:@917.4]
  wire  _T_36; // @[Lookup.scala 9:38:@919.4]
  wire  _T_40; // @[Lookup.scala 9:38:@921.4]
  wire [127:0] _T_43; // @[Lookup.scala 9:38:@922.4]
  wire  _T_44; // @[Lookup.scala 9:38:@923.4]
  wire  _T_48; // @[Lookup.scala 9:38:@925.4]
  wire  _T_52; // @[Lookup.scala 9:38:@927.4]
  wire  _T_56; // @[Lookup.scala 9:38:@929.4]
  wire  _T_58; // @[Lookup.scala 11:37:@931.4]
  wire  _T_59; // @[Lookup.scala 11:37:@932.4]
  wire  _T_60; // @[Lookup.scala 11:37:@933.4]
  wire  _T_61; // @[Lookup.scala 11:37:@934.4]
  wire  _T_62; // @[Lookup.scala 11:37:@935.4]
  wire  _T_63; // @[Lookup.scala 11:37:@936.4]
  wire  _T_64; // @[Lookup.scala 11:37:@937.4]
  wire  _T_65; // @[Lookup.scala 11:37:@938.4]
  wire  _T_66; // @[Lookup.scala 11:37:@939.4]
  wire  cs_val_inst; // @[Lookup.scala 11:37:@940.4]
  wire [2:0] _T_67; // @[Lookup.scala 11:37:@941.4]
  wire [2:0] _T_68; // @[Lookup.scala 11:37:@942.4]
  wire [2:0] _T_69; // @[Lookup.scala 11:37:@943.4]
  wire [2:0] _T_70; // @[Lookup.scala 11:37:@944.4]
  wire [2:0] _T_71; // @[Lookup.scala 11:37:@945.4]
  wire [2:0] _T_72; // @[Lookup.scala 11:37:@946.4]
  wire [2:0] _T_73; // @[Lookup.scala 11:37:@947.4]
  wire [2:0] _T_74; // @[Lookup.scala 11:37:@948.4]
  wire [2:0] _T_75; // @[Lookup.scala 11:37:@949.4]
  wire [2:0] _T_76; // @[Lookup.scala 11:37:@950.4]
  wire [2:0] cs_op_type; // @[Lookup.scala 11:37:@951.4]
  wire  _T_77; // @[Decode.scala 156:41:@952.4]
  wire  _T_79; // @[Decode.scala 157:44:@955.4]
  wire  _T_81; // @[Decode.scala 158:42:@958.4]
  assign _T_15 = io_inst & 128'h187; // @[Lookup.scala 9:38:@908.4]
  assign _T_16 = 128'h0 == _T_15; // @[Lookup.scala 9:38:@909.4]
  assign _T_20 = 128'h80 == _T_15; // @[Lookup.scala 9:38:@911.4]
  assign _T_24 = 128'h100 == _T_15; // @[Lookup.scala 9:38:@913.4]
  assign _T_28 = 128'h180 == _T_15; // @[Lookup.scala 9:38:@915.4]
  assign _T_31 = io_inst & 128'h7; // @[Lookup.scala 9:38:@916.4]
  assign _T_32 = 128'h1 == _T_31; // @[Lookup.scala 9:38:@917.4]
  assign _T_36 = 128'h2 == _T_31; // @[Lookup.scala 9:38:@919.4]
  assign _T_40 = 128'h3 == _T_31; // @[Lookup.scala 9:38:@921.4]
  assign _T_43 = io_inst & 128'h3000000000000000000000000007; // @[Lookup.scala 9:38:@922.4]
  assign _T_44 = 128'h4 == _T_43; // @[Lookup.scala 9:38:@923.4]
  assign _T_48 = 128'h1000000000000000000000000004 == _T_43; // @[Lookup.scala 9:38:@925.4]
  assign _T_52 = 128'h2000000000000000000000000004 == _T_43; // @[Lookup.scala 9:38:@927.4]
  assign _T_56 = 128'h3000000000000000000000000004 == _T_43; // @[Lookup.scala 9:38:@929.4]
  assign _T_58 = _T_52 ? 1'h1 : _T_56; // @[Lookup.scala 11:37:@931.4]
  assign _T_59 = _T_48 ? 1'h1 : _T_58; // @[Lookup.scala 11:37:@932.4]
  assign _T_60 = _T_44 ? 1'h1 : _T_59; // @[Lookup.scala 11:37:@933.4]
  assign _T_61 = _T_40 ? 1'h1 : _T_60; // @[Lookup.scala 11:37:@934.4]
  assign _T_62 = _T_36 ? 1'h1 : _T_61; // @[Lookup.scala 11:37:@935.4]
  assign _T_63 = _T_32 ? 1'h1 : _T_62; // @[Lookup.scala 11:37:@936.4]
  assign _T_64 = _T_28 ? 1'h1 : _T_63; // @[Lookup.scala 11:37:@937.4]
  assign _T_65 = _T_24 ? 1'h1 : _T_64; // @[Lookup.scala 11:37:@938.4]
  assign _T_66 = _T_20 ? 1'h1 : _T_65; // @[Lookup.scala 11:37:@939.4]
  assign cs_val_inst = _T_16 ? 1'h1 : _T_66; // @[Lookup.scala 11:37:@940.4]
  assign _T_67 = _T_56 ? 3'h2 : 3'h5; // @[Lookup.scala 11:37:@941.4]
  assign _T_68 = _T_52 ? 3'h2 : _T_67; // @[Lookup.scala 11:37:@942.4]
  assign _T_69 = _T_48 ? 3'h2 : _T_68; // @[Lookup.scala 11:37:@943.4]
  assign _T_70 = _T_44 ? 3'h2 : _T_69; // @[Lookup.scala 11:37:@944.4]
  assign _T_71 = _T_40 ? 3'h2 : _T_70; // @[Lookup.scala 11:37:@945.4]
  assign _T_72 = _T_36 ? 3'h2 : _T_71; // @[Lookup.scala 11:37:@946.4]
  assign _T_73 = _T_32 ? 3'h1 : _T_72; // @[Lookup.scala 11:37:@947.4]
  assign _T_74 = _T_28 ? 3'h2 : _T_73; // @[Lookup.scala 11:37:@948.4]
  assign _T_75 = _T_24 ? 3'h0 : _T_74; // @[Lookup.scala 11:37:@949.4]
  assign _T_76 = _T_20 ? 3'h0 : _T_75; // @[Lookup.scala 11:37:@950.4]
  assign cs_op_type = _T_16 ? 3'h2 : _T_76; // @[Lookup.scala 11:37:@951.4]
  assign _T_77 = cs_op_type == 3'h0; // @[Decode.scala 156:41:@952.4]
  assign _T_79 = cs_op_type == 3'h2; // @[Decode.scala 157:44:@955.4]
  assign _T_81 = cs_op_type == 3'h1; // @[Decode.scala 158:42:@958.4]
  assign io_isLoad = cs_val_inst & _T_77; // @[Decode.scala 156:13:@954.4]
  assign io_isCompute = cs_val_inst & _T_79; // @[Decode.scala 157:16:@957.4]
  assign io_isStore = cs_val_inst & _T_81; // @[Decode.scala 158:14:@960.4]
endmodule
module Fetch( // @[:@962.2]
  input          clock, // @[:@963.4]
  input          reset, // @[:@964.4]
  input          io_launch, // @[:@965.4]
  input  [31:0]  io_ins_baddr, // @[:@965.4]
  input  [31:0]  io_ins_count, // @[:@965.4]
  input          io_vme_rd_cmd_ready, // @[:@965.4]
  output         io_vme_rd_cmd_valid, // @[:@965.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@965.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@965.4]
  output         io_vme_rd_data_ready, // @[:@965.4]
  input          io_vme_rd_data_valid, // @[:@965.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@965.4]
  input          io_inst_ld_ready, // @[:@965.4]
  output         io_inst_ld_valid, // @[:@965.4]
  output [127:0] io_inst_ld_bits, // @[:@965.4]
  input          io_inst_co_ready, // @[:@965.4]
  output         io_inst_co_valid, // @[:@965.4]
  output [127:0] io_inst_co_bits, // @[:@965.4]
  input          io_inst_st_ready, // @[:@965.4]
  output         io_inst_st_valid, // @[:@965.4]
  output [127:0] io_inst_st_bits // @[:@965.4]
);
  wire  inst_q_clock; // @[Fetch.scala 57:22:@967.4]
  wire  inst_q_reset; // @[Fetch.scala 57:22:@967.4]
  wire  inst_q_io_enq_ready; // @[Fetch.scala 57:22:@967.4]
  wire  inst_q_io_enq_valid; // @[Fetch.scala 57:22:@967.4]
  wire [127:0] inst_q_io_enq_bits; // @[Fetch.scala 57:22:@967.4]
  wire  inst_q_io_deq_ready; // @[Fetch.scala 57:22:@967.4]
  wire  inst_q_io_deq_valid; // @[Fetch.scala 57:22:@967.4]
  wire [127:0] inst_q_io_deq_bits; // @[Fetch.scala 57:22:@967.4]
  wire [7:0] inst_q_io_count; // @[Fetch.scala 57:22:@967.4]
  wire [127:0] dec_io_inst; // @[Fetch.scala 58:19:@970.4]
  wire  dec_io_isLoad; // @[Fetch.scala 58:19:@970.4]
  wire  dec_io_isCompute; // @[Fetch.scala 58:19:@970.4]
  wire  dec_io_isStore; // @[Fetch.scala 58:19:@970.4]
  reg  s1_launch; // @[Fetch.scala 60:26:@973.4]
  reg [31:0] _RAND_0;
  wire  _T_65; // @[Fetch.scala 61:27:@975.4]
  wire  pulse; // @[Fetch.scala 61:25:@976.4]
  reg [31:0] raddr; // @[Fetch.scala 63:18:@977.4]
  reg [31:0] _RAND_1;
  reg [7:0] rlen; // @[Fetch.scala 64:17:@978.4]
  reg [31:0] _RAND_2;
  reg [7:0] ilen; // @[Fetch.scala 65:17:@979.4]
  reg [31:0] _RAND_3;
  reg [31:0] xrem; // @[Fetch.scala 67:17:@980.4]
  reg [31:0] _RAND_4;
  wire [32:0] _GEN_46; // @[Fetch.scala 68:29:@981.4]
  wire [32:0] _T_71; // @[Fetch.scala 68:29:@981.4]
  wire [33:0] _T_73; // @[Fetch.scala 68:37:@982.4]
  wire [33:0] _T_74; // @[Fetch.scala 68:37:@983.4]
  wire [32:0] xsize; // @[Fetch.scala 68:37:@984.4]
  reg [2:0] state; // @[Fetch.scala 73:22:@985.4]
  reg [31:0] _RAND_5;
  wire  _T_76; // @[Conditional.scala 37:30:@986.4]
  wire  _T_77; // @[Fetch.scala 80:20:@990.8]
  wire [32:0] _T_79; // @[Fetch.scala 82:25:@993.10]
  wire [9:0] _T_82; // @[Fetch.scala 85:24:@998.10]
  wire [9:0] _T_83; // @[Fetch.scala 85:24:@999.10]
  wire [8:0] _T_84; // @[Fetch.scala 85:24:@1000.10]
  wire [8:0] _T_86; // @[Fetch.scala 86:25:@1002.10]
  wire [9:0] _T_88; // @[Fetch.scala 86:33:@1003.10]
  wire [9:0] _T_89; // @[Fetch.scala 86:33:@1004.10]
  wire [8:0] _T_90; // @[Fetch.scala 86:33:@1005.10]
  wire [33:0] _T_91; // @[Fetch.scala 87:25:@1007.10]
  wire [33:0] _T_92; // @[Fetch.scala 87:25:@1008.10]
  wire [32:0] _T_93; // @[Fetch.scala 87:25:@1009.10]
  wire [32:0] _GEN_0; // @[Fetch.scala 80:28:@991.8]
  wire [32:0] _GEN_1; // @[Fetch.scala 80:28:@991.8]
  wire [32:0] _GEN_2; // @[Fetch.scala 80:28:@991.8]
  wire [2:0] _GEN_3; // @[Fetch.scala 78:19:@988.6]
  wire [32:0] _GEN_4; // @[Fetch.scala 78:19:@988.6]
  wire [32:0] _GEN_5; // @[Fetch.scala 78:19:@988.6]
  wire [32:0] _GEN_6; // @[Fetch.scala 78:19:@988.6]
  wire  _T_94; // @[Conditional.scala 37:30:@1015.6]
  wire [2:0] _GEN_7; // @[Fetch.scala 92:33:@1017.8]
  wire  _T_95; // @[Conditional.scala 37:30:@1022.8]
  wire [2:0] _GEN_8; // @[Fetch.scala 97:34:@1024.10]
  wire  _T_96; // @[Conditional.scala 37:30:@1029.10]
  wire  _T_97; // @[Fetch.scala 103:30:@1032.14]
  wire [2:0] _GEN_9; // @[Fetch.scala 103:40:@1033.14]
  wire [2:0] _GEN_10; // @[Fetch.scala 102:34:@1031.12]
  wire  _T_98; // @[Conditional.scala 37:30:@1042.12]
  wire  _T_100; // @[Fetch.scala 111:28:@1044.14]
  wire  _T_102; // @[Fetch.scala 112:19:@1046.16]
  wire  _T_103; // @[Fetch.scala 114:25:@1051.18]
  wire [31:0] _T_105; // @[Fetch.scala 117:24:@1055.20]
  wire [32:0] _T_117; // @[Fetch.scala 123:24:@1070.20]
  wire [32:0] _T_118; // @[Fetch.scala 123:24:@1071.20]
  wire [31:0] _T_119; // @[Fetch.scala 123:24:@1072.20]
  wire [31:0] _GEN_12; // @[Fetch.scala 114:33:@1052.18]
  wire [31:0] _GEN_13; // @[Fetch.scala 114:33:@1052.18]
  wire [31:0] _GEN_14; // @[Fetch.scala 114:33:@1052.18]
  wire [2:0] _GEN_15; // @[Fetch.scala 112:28:@1047.16]
  wire [31:0] _GEN_16; // @[Fetch.scala 112:28:@1047.16]
  wire [31:0] _GEN_17; // @[Fetch.scala 112:28:@1047.16]
  wire [31:0] _GEN_18; // @[Fetch.scala 112:28:@1047.16]
  wire [2:0] _GEN_19; // @[Fetch.scala 111:37:@1045.14]
  wire [31:0] _GEN_20; // @[Fetch.scala 111:37:@1045.14]
  wire [31:0] _GEN_21; // @[Fetch.scala 111:37:@1045.14]
  wire [31:0] _GEN_22; // @[Fetch.scala 111:37:@1045.14]
  wire [2:0] _GEN_23; // @[Conditional.scala 39:67:@1043.12]
  wire [31:0] _GEN_24; // @[Conditional.scala 39:67:@1043.12]
  wire [31:0] _GEN_25; // @[Conditional.scala 39:67:@1043.12]
  wire [31:0] _GEN_26; // @[Conditional.scala 39:67:@1043.12]
  wire [2:0] _GEN_27; // @[Conditional.scala 39:67:@1030.10]
  wire [31:0] _GEN_28; // @[Conditional.scala 39:67:@1030.10]
  wire [31:0] _GEN_29; // @[Conditional.scala 39:67:@1030.10]
  wire [31:0] _GEN_30; // @[Conditional.scala 39:67:@1030.10]
  wire [2:0] _GEN_31; // @[Conditional.scala 39:67:@1023.8]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67:@1023.8]
  wire [31:0] _GEN_33; // @[Conditional.scala 39:67:@1023.8]
  wire [31:0] _GEN_34; // @[Conditional.scala 39:67:@1023.8]
  wire [2:0] _GEN_35; // @[Conditional.scala 39:67:@1016.6]
  wire [31:0] _GEN_36; // @[Conditional.scala 39:67:@1016.6]
  wire [31:0] _GEN_37; // @[Conditional.scala 39:67:@1016.6]
  wire [31:0] _GEN_38; // @[Conditional.scala 39:67:@1016.6]
  wire [2:0] _GEN_39; // @[Conditional.scala 40:58:@987.4]
  wire [32:0] _GEN_40; // @[Conditional.scala 40:58:@987.4]
  wire [32:0] _GEN_41; // @[Conditional.scala 40:58:@987.4]
  wire [32:0] _GEN_42; // @[Conditional.scala 40:58:@987.4]
  wire  _T_120; // @[Fetch.scala 130:14:@1077.4]
  wire  _T_121; // @[Fetch.scala 132:20:@1082.6]
  wire  _T_124; // @[Fetch.scala 132:31:@1084.6]
  wire  _T_126; // @[Fetch.scala 132:66:@1085.6]
  wire  _T_127; // @[Fetch.scala 132:58:@1086.6]
  wire [32:0] _T_128; // @[Fetch.scala 133:20:@1088.8]
  wire [31:0] _T_129; // @[Fetch.scala 133:20:@1089.8]
  wire [31:0] _GEN_43; // @[Fetch.scala 132:75:@1087.6]
  reg [63:0] lsb; // @[Fetch.scala 142:16:@1097.4]
  reg [63:0] _RAND_6;
  wire  _T_132; // @[Fetch.scala 146:14:@1099.4]
  wire  _T_133; // @[Fetch.scala 148:55:@1103.4]
  wire  _T_135; // @[Fetch.scala 155:37:@1108.4]
  wire  _T_138; // @[Fetch.scala 156:40:@1112.4]
  wire  _T_141; // @[Fetch.scala 157:38:@1116.4]
  wire [2:0] deq_sel; // @[Cat.scala 30:58:@1124.4]
  wire  _T_149; // @[Mux.scala 46:19:@1125.4]
  wire  _T_150; // @[Mux.scala 46:16:@1126.4]
  wire  _T_151; // @[Mux.scala 46:19:@1127.4]
  wire  _T_152; // @[Mux.scala 46:16:@1128.4]
  wire  _T_153; // @[Mux.scala 46:19:@1129.4]
  wire  deq_ready; // @[Mux.scala 46:16:@1130.4]
  wire  _T_154; // @[Fetch.scala 175:36:@1131.4]
  Queue inst_q ( // @[Fetch.scala 57:22:@967.4]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits),
    .io_count(inst_q_io_count)
  );
  FetchDecode dec ( // @[Fetch.scala 58:19:@970.4]
    .io_inst(dec_io_inst),
    .io_isLoad(dec_io_isLoad),
    .io_isCompute(dec_io_isCompute),
    .io_isStore(dec_io_isStore)
  );
  assign _T_65 = ~ s1_launch; // @[Fetch.scala 61:27:@975.4]
  assign pulse = io_launch & _T_65; // @[Fetch.scala 61:25:@976.4]
  assign _GEN_46 = {{1'd0}, io_ins_count}; // @[Fetch.scala 68:29:@981.4]
  assign _T_71 = _GEN_46 << 1'h1; // @[Fetch.scala 68:29:@981.4]
  assign _T_73 = _T_71 - 33'h1; // @[Fetch.scala 68:37:@982.4]
  assign _T_74 = $unsigned(_T_73); // @[Fetch.scala 68:37:@983.4]
  assign xsize = _T_74[32:0]; // @[Fetch.scala 68:37:@984.4]
  assign _T_76 = 3'h0 == state; // @[Conditional.scala 37:30:@986.4]
  assign _T_77 = xsize < 33'h100; // @[Fetch.scala 80:20:@990.8]
  assign _T_79 = xsize >> 1'h1; // @[Fetch.scala 82:25:@993.10]
  assign _T_82 = 9'h100 - 9'h1; // @[Fetch.scala 85:24:@998.10]
  assign _T_83 = $unsigned(_T_82); // @[Fetch.scala 85:24:@999.10]
  assign _T_84 = _T_83[8:0]; // @[Fetch.scala 85:24:@1000.10]
  assign _T_86 = 9'h100 >> 1'h1; // @[Fetch.scala 86:25:@1002.10]
  assign _T_88 = _T_86 - 9'h1; // @[Fetch.scala 86:33:@1003.10]
  assign _T_89 = $unsigned(_T_88); // @[Fetch.scala 86:33:@1004.10]
  assign _T_90 = _T_89[8:0]; // @[Fetch.scala 86:33:@1005.10]
  assign _T_91 = xsize - 33'h100; // @[Fetch.scala 87:25:@1007.10]
  assign _T_92 = $unsigned(_T_91); // @[Fetch.scala 87:25:@1008.10]
  assign _T_93 = _T_92[32:0]; // @[Fetch.scala 87:25:@1009.10]
  assign _GEN_0 = _T_77 ? xsize : {{24'd0}, _T_84}; // @[Fetch.scala 80:28:@991.8]
  assign _GEN_1 = _T_77 ? _T_79 : {{24'd0}, _T_90}; // @[Fetch.scala 80:28:@991.8]
  assign _GEN_2 = _T_77 ? 33'h0 : _T_93; // @[Fetch.scala 80:28:@991.8]
  assign _GEN_3 = pulse ? 3'h1 : state; // @[Fetch.scala 78:19:@988.6]
  assign _GEN_4 = pulse ? _GEN_0 : {{25'd0}, rlen}; // @[Fetch.scala 78:19:@988.6]
  assign _GEN_5 = pulse ? _GEN_1 : {{25'd0}, ilen}; // @[Fetch.scala 78:19:@988.6]
  assign _GEN_6 = pulse ? _GEN_2 : {{1'd0}, xrem}; // @[Fetch.scala 78:19:@988.6]
  assign _T_94 = 3'h1 == state; // @[Conditional.scala 37:30:@1015.6]
  assign _GEN_7 = io_vme_rd_cmd_ready ? 3'h2 : state; // @[Fetch.scala 92:33:@1017.8]
  assign _T_95 = 3'h2 == state; // @[Conditional.scala 37:30:@1022.8]
  assign _GEN_8 = io_vme_rd_data_valid ? 3'h3 : state; // @[Fetch.scala 97:34:@1024.10]
  assign _T_96 = 3'h3 == state; // @[Conditional.scala 37:30:@1029.10]
  assign _T_97 = inst_q_io_count == ilen; // @[Fetch.scala 103:30:@1032.14]
  assign _GEN_9 = _T_97 ? 3'h4 : 3'h2; // @[Fetch.scala 103:40:@1033.14]
  assign _GEN_10 = io_vme_rd_data_valid ? _GEN_9 : state; // @[Fetch.scala 102:34:@1031.12]
  assign _T_98 = 3'h4 == state; // @[Conditional.scala 37:30:@1042.12]
  assign _T_100 = inst_q_io_count == 8'h0; // @[Fetch.scala 111:28:@1044.14]
  assign _T_102 = xrem == 32'h0; // @[Fetch.scala 112:19:@1046.16]
  assign _T_103 = xrem < 32'h100; // @[Fetch.scala 114:25:@1051.18]
  assign _T_105 = xrem >> 1'h1; // @[Fetch.scala 117:24:@1055.20]
  assign _T_117 = xrem - 32'h100; // @[Fetch.scala 123:24:@1070.20]
  assign _T_118 = $unsigned(_T_117); // @[Fetch.scala 123:24:@1071.20]
  assign _T_119 = _T_118[31:0]; // @[Fetch.scala 123:24:@1072.20]
  assign _GEN_12 = _T_103 ? xrem : {{23'd0}, _T_84}; // @[Fetch.scala 114:33:@1052.18]
  assign _GEN_13 = _T_103 ? _T_105 : {{23'd0}, _T_90}; // @[Fetch.scala 114:33:@1052.18]
  assign _GEN_14 = _T_103 ? 32'h0 : _T_119; // @[Fetch.scala 114:33:@1052.18]
  assign _GEN_15 = _T_102 ? 3'h0 : 3'h1; // @[Fetch.scala 112:28:@1047.16]
  assign _GEN_16 = _T_102 ? {{24'd0}, rlen} : _GEN_12; // @[Fetch.scala 112:28:@1047.16]
  assign _GEN_17 = _T_102 ? {{24'd0}, ilen} : _GEN_13; // @[Fetch.scala 112:28:@1047.16]
  assign _GEN_18 = _T_102 ? xrem : _GEN_14; // @[Fetch.scala 112:28:@1047.16]
  assign _GEN_19 = _T_100 ? _GEN_15 : state; // @[Fetch.scala 111:37:@1045.14]
  assign _GEN_20 = _T_100 ? _GEN_16 : {{24'd0}, rlen}; // @[Fetch.scala 111:37:@1045.14]
  assign _GEN_21 = _T_100 ? _GEN_17 : {{24'd0}, ilen}; // @[Fetch.scala 111:37:@1045.14]
  assign _GEN_22 = _T_100 ? _GEN_18 : xrem; // @[Fetch.scala 111:37:@1045.14]
  assign _GEN_23 = _T_98 ? _GEN_19 : state; // @[Conditional.scala 39:67:@1043.12]
  assign _GEN_24 = _T_98 ? _GEN_20 : {{24'd0}, rlen}; // @[Conditional.scala 39:67:@1043.12]
  assign _GEN_25 = _T_98 ? _GEN_21 : {{24'd0}, ilen}; // @[Conditional.scala 39:67:@1043.12]
  assign _GEN_26 = _T_98 ? _GEN_22 : xrem; // @[Conditional.scala 39:67:@1043.12]
  assign _GEN_27 = _T_96 ? _GEN_10 : _GEN_23; // @[Conditional.scala 39:67:@1030.10]
  assign _GEN_28 = _T_96 ? {{24'd0}, rlen} : _GEN_24; // @[Conditional.scala 39:67:@1030.10]
  assign _GEN_29 = _T_96 ? {{24'd0}, ilen} : _GEN_25; // @[Conditional.scala 39:67:@1030.10]
  assign _GEN_30 = _T_96 ? xrem : _GEN_26; // @[Conditional.scala 39:67:@1030.10]
  assign _GEN_31 = _T_95 ? _GEN_8 : _GEN_27; // @[Conditional.scala 39:67:@1023.8]
  assign _GEN_32 = _T_95 ? {{24'd0}, rlen} : _GEN_28; // @[Conditional.scala 39:67:@1023.8]
  assign _GEN_33 = _T_95 ? {{24'd0}, ilen} : _GEN_29; // @[Conditional.scala 39:67:@1023.8]
  assign _GEN_34 = _T_95 ? xrem : _GEN_30; // @[Conditional.scala 39:67:@1023.8]
  assign _GEN_35 = _T_94 ? _GEN_7 : _GEN_31; // @[Conditional.scala 39:67:@1016.6]
  assign _GEN_36 = _T_94 ? {{24'd0}, rlen} : _GEN_32; // @[Conditional.scala 39:67:@1016.6]
  assign _GEN_37 = _T_94 ? {{24'd0}, ilen} : _GEN_33; // @[Conditional.scala 39:67:@1016.6]
  assign _GEN_38 = _T_94 ? xrem : _GEN_34; // @[Conditional.scala 39:67:@1016.6]
  assign _GEN_39 = _T_76 ? _GEN_3 : _GEN_35; // @[Conditional.scala 40:58:@987.4]
  assign _GEN_40 = _T_76 ? _GEN_4 : {{1'd0}, _GEN_36}; // @[Conditional.scala 40:58:@987.4]
  assign _GEN_41 = _T_76 ? _GEN_5 : {{1'd0}, _GEN_37}; // @[Conditional.scala 40:58:@987.4]
  assign _GEN_42 = _T_76 ? _GEN_6 : {{1'd0}, _GEN_38}; // @[Conditional.scala 40:58:@987.4]
  assign _T_120 = state == 3'h0; // @[Fetch.scala 130:14:@1077.4]
  assign _T_121 = state == 3'h4; // @[Fetch.scala 132:20:@1082.6]
  assign _T_124 = _T_121 & _T_100; // @[Fetch.scala 132:31:@1084.6]
  assign _T_126 = xrem != 32'h0; // @[Fetch.scala 132:66:@1085.6]
  assign _T_127 = _T_124 & _T_126; // @[Fetch.scala 132:58:@1086.6]
  assign _T_128 = raddr + 32'h800; // @[Fetch.scala 133:20:@1088.8]
  assign _T_129 = raddr + 32'h800; // @[Fetch.scala 133:20:@1089.8]
  assign _GEN_43 = _T_127 ? _T_129 : raddr; // @[Fetch.scala 132:75:@1087.6]
  assign _T_132 = state == 3'h2; // @[Fetch.scala 146:14:@1099.4]
  assign _T_133 = state == 3'h3; // @[Fetch.scala 148:55:@1103.4]
  assign _T_135 = dec_io_isLoad & inst_q_io_deq_valid; // @[Fetch.scala 155:37:@1108.4]
  assign _T_138 = dec_io_isCompute & inst_q_io_deq_valid; // @[Fetch.scala 156:40:@1112.4]
  assign _T_141 = dec_io_isStore & inst_q_io_deq_valid; // @[Fetch.scala 157:38:@1116.4]
  assign deq_sel = {dec_io_isCompute,dec_io_isStore,dec_io_isLoad}; // @[Cat.scala 30:58:@1124.4]
  assign _T_149 = 3'h4 == deq_sel; // @[Mux.scala 46:19:@1125.4]
  assign _T_150 = _T_149 ? io_inst_co_ready : 1'h0; // @[Mux.scala 46:16:@1126.4]
  assign _T_151 = 3'h2 == deq_sel; // @[Mux.scala 46:19:@1127.4]
  assign _T_152 = _T_151 ? io_inst_st_ready : _T_150; // @[Mux.scala 46:16:@1128.4]
  assign _T_153 = 3'h1 == deq_sel; // @[Mux.scala 46:19:@1129.4]
  assign deq_ready = _T_153 ? io_inst_ld_ready : _T_152; // @[Mux.scala 46:16:@1130.4]
  assign _T_154 = deq_ready & inst_q_io_deq_valid; // @[Fetch.scala 175:36:@1131.4]
  assign io_vme_rd_cmd_valid = state == 3'h1; // @[Fetch.scala 136:23:@1093.4]
  assign io_vme_rd_cmd_bits_addr = raddr; // @[Fetch.scala 137:27:@1094.4]
  assign io_vme_rd_cmd_bits_len = rlen; // @[Fetch.scala 138:26:@1095.4]
  assign io_vme_rd_data_ready = inst_q_io_enq_ready; // @[Fetch.scala 140:24:@1096.4]
  assign io_inst_ld_valid = _T_135 & _T_121; // @[Fetch.scala 155:20:@1111.4]
  assign io_inst_ld_bits = inst_q_io_deq_bits; // @[Fetch.scala 159:19:@1120.4]
  assign io_inst_co_valid = _T_138 & _T_121; // @[Fetch.scala 156:20:@1115.4]
  assign io_inst_co_bits = inst_q_io_deq_bits; // @[Fetch.scala 160:19:@1121.4]
  assign io_inst_st_valid = _T_141 & _T_121; // @[Fetch.scala 157:20:@1119.4]
  assign io_inst_st_bits = inst_q_io_deq_bits; // @[Fetch.scala 161:19:@1122.4]
  assign inst_q_clock = clock; // @[:@968.4]
  assign inst_q_reset = reset; // @[:@969.4]
  assign inst_q_io_enq_valid = io_vme_rd_data_valid & _T_133; // @[Fetch.scala 148:23:@1105.4]
  assign inst_q_io_enq_bits = {io_vme_rd_data_bits,lsb}; // @[Fetch.scala 149:22:@1106.4]
  assign inst_q_io_deq_ready = _T_154 & _T_121; // @[Fetch.scala 175:23:@1134.4]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Fetch.scala 152:15:@1107.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_launch = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  raddr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rlen = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ilen = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xrem = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{`RANDOM}};
  lsb = _RAND_6[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    s1_launch <= io_launch;
    if (_T_120) begin
      raddr <= io_ins_baddr;
    end else begin
      if (_T_127) begin
        raddr <= _T_129;
      end
    end
    rlen <= _GEN_40[7:0];
    ilen <= _GEN_41[7:0];
    xrem <= _GEN_42[31:0];
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_76) begin
        if (pulse) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_94) begin
          if (io_vme_rd_cmd_ready) begin
            state <= 3'h2;
          end
        end else begin
          if (_T_95) begin
            if (io_vme_rd_data_valid) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_96) begin
              if (io_vme_rd_data_valid) begin
                if (_T_97) begin
                  state <= 3'h4;
                end else begin
                  state <= 3'h2;
                end
              end
            end else begin
              if (_T_98) begin
                if (_T_100) begin
                  if (_T_102) begin
                    state <= 3'h0;
                  end else begin
                    state <= 3'h1;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_132) begin
      lsb <= io_vme_rd_data_bits;
    end
  end
endmodule
module Semaphore( // @[:@1136.2]
  input   clock, // @[:@1137.4]
  input   reset, // @[:@1138.4]
  input   io_spost, // @[:@1139.4]
  input   io_swait, // @[:@1139.4]
  output  io_sready // @[:@1139.4]
);
  reg [7:0] cnt; // @[Semaphore.scala 38:20:@1141.4]
  reg [31:0] _RAND_0;
  wire  _T_14; // @[Semaphore.scala 39:20:@1142.4]
  wire  _T_15; // @[Semaphore.scala 39:17:@1143.4]
  wire  _T_17; // @[Semaphore.scala 39:37:@1144.4]
  wire  _T_18; // @[Semaphore.scala 39:30:@1145.4]
  wire [8:0] _T_20; // @[Semaphore.scala 40:16:@1147.6]
  wire [7:0] _T_21; // @[Semaphore.scala 40:16:@1148.6]
  wire [7:0] _GEN_0; // @[Semaphore.scala 39:74:@1146.4]
  wire  _T_23; // @[Semaphore.scala 42:8:@1151.4]
  wire  _T_24; // @[Semaphore.scala 42:18:@1152.4]
  wire  _T_26; // @[Semaphore.scala 42:37:@1153.4]
  wire  _T_27; // @[Semaphore.scala 42:30:@1154.4]
  wire [8:0] _T_29; // @[Semaphore.scala 42:59:@1156.6]
  wire [8:0] _T_30; // @[Semaphore.scala 42:59:@1157.6]
  wire [7:0] _T_31; // @[Semaphore.scala 42:59:@1158.6]
  wire [7:0] _GEN_1; // @[Semaphore.scala 42:46:@1155.4]
  assign _T_14 = io_swait == 1'h0; // @[Semaphore.scala 39:20:@1142.4]
  assign _T_15 = io_spost & _T_14; // @[Semaphore.scala 39:17:@1143.4]
  assign _T_17 = cnt != 8'hff; // @[Semaphore.scala 39:37:@1144.4]
  assign _T_18 = _T_15 & _T_17; // @[Semaphore.scala 39:30:@1145.4]
  assign _T_20 = cnt + 8'h1; // @[Semaphore.scala 40:16:@1147.6]
  assign _T_21 = cnt + 8'h1; // @[Semaphore.scala 40:16:@1148.6]
  assign _GEN_0 = _T_18 ? _T_21 : cnt; // @[Semaphore.scala 39:74:@1146.4]
  assign _T_23 = io_spost == 1'h0; // @[Semaphore.scala 42:8:@1151.4]
  assign _T_24 = _T_23 & io_swait; // @[Semaphore.scala 42:18:@1152.4]
  assign _T_26 = cnt != 8'h0; // @[Semaphore.scala 42:37:@1153.4]
  assign _T_27 = _T_24 & _T_26; // @[Semaphore.scala 42:30:@1154.4]
  assign _T_29 = cnt - 8'h1; // @[Semaphore.scala 42:59:@1156.6]
  assign _T_30 = $unsigned(_T_29); // @[Semaphore.scala 42:59:@1157.6]
  assign _T_31 = _T_30[7:0]; // @[Semaphore.scala 42:59:@1158.6]
  assign _GEN_1 = _T_27 ? _T_31 : _GEN_0; // @[Semaphore.scala 42:46:@1155.4]
  assign io_sready = cnt != 8'h0; // @[Semaphore.scala 43:13:@1162.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 8'h0;
    end else begin
      if (_T_27) begin
        cnt <= _T_31;
      end else begin
        if (_T_18) begin
          cnt <= _T_21;
        end
      end
    end
  end
endmodule
module Queue_1( // @[:@1164.2]
  input          clock, // @[:@1165.4]
  input          reset, // @[:@1166.4]
  output         io_enq_ready, // @[:@1167.4]
  input          io_enq_valid, // @[:@1167.4]
  input  [127:0] io_enq_bits, // @[:@1167.4]
  input          io_deq_ready, // @[:@1167.4]
  output         io_deq_valid, // @[:@1167.4]
  output [127:0] io_deq_bits // @[:@1167.4]
);
  reg [127:0] _T_35 [0:511]; // @[Decoupled.scala 215:24:@1169.4]
  reg [127:0] _RAND_0;
  wire [127:0] _T_35__T_68_data; // @[Decoupled.scala 215:24:@1169.4]
  wire [8:0] _T_35__T_68_addr; // @[Decoupled.scala 215:24:@1169.4]
  wire [127:0] _T_35__T_54_data; // @[Decoupled.scala 215:24:@1169.4]
  wire [8:0] _T_35__T_54_addr; // @[Decoupled.scala 215:24:@1169.4]
  wire  _T_35__T_54_mask; // @[Decoupled.scala 215:24:@1169.4]
  wire  _T_35__T_54_en; // @[Decoupled.scala 215:24:@1169.4]
  reg [8:0] value; // @[Counter.scala 26:33:@1170.4]
  reg [31:0] _RAND_1;
  reg [8:0] value_1; // @[Counter.scala 26:33:@1171.4]
  reg [31:0] _RAND_2;
  reg  _T_42; // @[Decoupled.scala 218:35:@1172.4]
  reg [31:0] _RAND_3;
  wire  _T_43; // @[Decoupled.scala 220:41:@1173.4]
  wire  _T_45; // @[Decoupled.scala 221:36:@1174.4]
  wire  _T_46; // @[Decoupled.scala 221:33:@1175.4]
  wire  _T_47; // @[Decoupled.scala 222:32:@1176.4]
  wire  _T_48; // @[Decoupled.scala 37:37:@1177.4]
  wire  _T_51; // @[Decoupled.scala 37:37:@1180.4]
  wire [9:0] _T_57; // @[Counter.scala 35:22:@1187.6]
  wire [8:0] _T_58; // @[Counter.scala 35:22:@1188.6]
  wire [8:0] _GEN_5; // @[Decoupled.scala 226:17:@1183.4]
  wire [9:0] _T_61; // @[Counter.scala 35:22:@1193.6]
  wire [8:0] _T_62; // @[Counter.scala 35:22:@1194.6]
  wire [8:0] _GEN_6; // @[Decoupled.scala 230:17:@1191.4]
  wire  _T_63; // @[Decoupled.scala 233:16:@1197.4]
  wire  _GEN_7; // @[Decoupled.scala 233:28:@1198.4]
  assign _T_35__T_68_addr = value_1;
  assign _T_35__T_68_data = _T_35[_T_35__T_68_addr]; // @[Decoupled.scala 215:24:@1169.4]
  assign _T_35__T_54_data = io_enq_bits;
  assign _T_35__T_54_addr = value;
  assign _T_35__T_54_mask = 1'h1;
  assign _T_35__T_54_en = io_enq_ready & io_enq_valid;
  assign _T_43 = value == value_1; // @[Decoupled.scala 220:41:@1173.4]
  assign _T_45 = _T_42 == 1'h0; // @[Decoupled.scala 221:36:@1174.4]
  assign _T_46 = _T_43 & _T_45; // @[Decoupled.scala 221:33:@1175.4]
  assign _T_47 = _T_43 & _T_42; // @[Decoupled.scala 222:32:@1176.4]
  assign _T_48 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37:@1177.4]
  assign _T_51 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37:@1180.4]
  assign _T_57 = value + 9'h1; // @[Counter.scala 35:22:@1187.6]
  assign _T_58 = value + 9'h1; // @[Counter.scala 35:22:@1188.6]
  assign _GEN_5 = _T_48 ? _T_58 : value; // @[Decoupled.scala 226:17:@1183.4]
  assign _T_61 = value_1 + 9'h1; // @[Counter.scala 35:22:@1193.6]
  assign _T_62 = value_1 + 9'h1; // @[Counter.scala 35:22:@1194.6]
  assign _GEN_6 = _T_51 ? _T_62 : value_1; // @[Decoupled.scala 230:17:@1191.4]
  assign _T_63 = _T_48 != _T_51; // @[Decoupled.scala 233:16:@1197.4]
  assign _GEN_7 = _T_63 ? _T_48 : _T_42; // @[Decoupled.scala 233:28:@1198.4]
  assign io_enq_ready = _T_47 == 1'h0; // @[Decoupled.scala 238:16:@1204.4]
  assign io_deq_valid = _T_46 == 1'h0; // @[Decoupled.scala 237:16:@1202.4]
  assign io_deq_bits = _T_35__T_68_data; // @[Decoupled.scala 239:15:@1206.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    _T_35[initvar] = _RAND_0[127:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_42 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_35__T_54_en & _T_35__T_54_mask) begin
      _T_35[_T_35__T_54_addr] <= _T_35__T_54_data; // @[Decoupled.scala 215:24:@1169.4]
    end
    if (reset) begin
      value <= 9'h0;
    end else begin
      if (_T_48) begin
        value <= _T_58;
      end
    end
    if (reset) begin
      value_1 <= 9'h0;
    end else begin
      if (_T_51) begin
        value_1 <= _T_62;
      end
    end
    if (reset) begin
      _T_42 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_42 <= _T_48;
      end
    end
  end
endmodule
module LoadDecode( // @[:@1215.2]
  input  [127:0] io_inst, // @[:@1218.4]
  output         io_push_next, // @[:@1218.4]
  output         io_pop_next, // @[:@1218.4]
  output         io_isInput, // @[:@1218.4]
  output         io_isWeight, // @[:@1218.4]
  output         io_isSync // @[:@1218.4]
);
  wire [15:0] dec_xsize; // @[Decode.scala 174:29:@1243.4]
  wire [127:0] _T_39; // @[Decode.scala 177:25:@1257.4]
  wire  _T_40; // @[Decode.scala 177:25:@1258.4]
  wire  _T_42; // @[Decode.scala 177:46:@1259.4]
  wire  _T_47; // @[Decode.scala 178:26:@1263.4]
  wire  _T_59; // @[Decode.scala 179:34:@1271.4]
  wire  _T_61; // @[Decode.scala 179:66:@1272.4]
  assign dec_xsize = io_inst[95:80]; // @[Decode.scala 174:29:@1243.4]
  assign _T_39 = io_inst & 128'h187; // @[Decode.scala 177:25:@1257.4]
  assign _T_40 = 128'h100 == _T_39; // @[Decode.scala 177:25:@1258.4]
  assign _T_42 = dec_xsize != 16'h0; // @[Decode.scala 177:46:@1259.4]
  assign _T_47 = 128'h80 == _T_39; // @[Decode.scala 178:26:@1263.4]
  assign _T_59 = _T_40 | _T_47; // @[Decode.scala 179:34:@1271.4]
  assign _T_61 = dec_xsize == 16'h0; // @[Decode.scala 179:66:@1272.4]
  assign io_push_next = io_inst[6]; // @[Decode.scala 175:16:@1255.4]
  assign io_pop_next = io_inst[4]; // @[Decode.scala 176:15:@1256.4]
  assign io_isInput = _T_40 & _T_42; // @[Decode.scala 177:14:@1261.4]
  assign io_isWeight = _T_47 & _T_42; // @[Decode.scala 178:15:@1266.4]
  assign io_isSync = _T_59 & _T_61; // @[Decode.scala 179:13:@1274.4]
endmodule
module TensorDataCtrl( // @[:@1276.2]
  input          clock, // @[:@1277.4]
  input          io_start, // @[:@1279.4]
  output         io_done, // @[:@1279.4]
  input  [127:0] io_inst, // @[:@1279.4]
  input  [31:0]  io_baddr, // @[:@1279.4]
  input          io_xinit, // @[:@1279.4]
  input          io_xupdate, // @[:@1279.4]
  input          io_yupdate, // @[:@1279.4]
  output         io_stride, // @[:@1279.4]
  output         io_split, // @[:@1279.4]
  output [31:0]  io_addr, // @[:@1279.4]
  output [7:0]   io_len // @[:@1279.4]
);
  wire [31:0] dec_dram_offset; // @[TensorUtil.scala 251:29:@1298.4]
  wire [15:0] dec_ysize; // @[TensorUtil.scala 251:29:@1302.4]
  wire [15:0] dec_xsize; // @[TensorUtil.scala 251:29:@1304.4]
  wire [15:0] dec_xstride; // @[TensorUtil.scala 251:29:@1306.4]
  reg [31:0] caddr; // @[TensorUtil.scala 253:18:@1316.4]
  reg [31:0] _RAND_0;
  reg [31:0] baddr; // @[TensorUtil.scala 254:18:@1317.4]
  reg [31:0] _RAND_1;
  reg [7:0] len; // @[TensorUtil.scala 255:16:@1318.4]
  reg [31:0] _RAND_2;
  reg [7:0] xcnt; // @[TensorUtil.scala 267:17:@1383.4]
  reg [31:0] _RAND_3;
  reg [15:0] xrem; // @[TensorUtil.scala 268:17:@1384.4]
  reg [31:0] _RAND_4;
  wire [16:0] _GEN_27; // @[TensorUtil.scala 269:26:@1385.4]
  wire [16:0] _T_154; // @[TensorUtil.scala 269:26:@1385.4]
  wire [17:0] _T_156; // @[TensorUtil.scala 269:51:@1386.4]
  wire [17:0] _T_157; // @[TensorUtil.scala 269:51:@1387.4]
  wire [16:0] xsize; // @[TensorUtil.scala 269:51:@1388.4]
  reg [15:0] ycnt; // @[TensorUtil.scala 271:17:@1389.4]
  reg [31:0] _RAND_5;
  reg [31:0] xfer_bytes; // @[TensorUtil.scala 273:23:@1390.4]
  reg [31:0] _RAND_6;
  wire [19:0] _GEN_28; // @[TensorUtil.scala 275:35:@1391.4]
  wire [19:0] xstride_bytes; // @[TensorUtil.scala 275:35:@1391.4]
  wire [35:0] _GEN_29; // @[TensorUtil.scala 277:66:@1392.4]
  wire [35:0] _T_160; // @[TensorUtil.scala 277:66:@1392.4]
  wire [35:0] _T_161; // @[TensorUtil.scala 277:47:@1393.4]
  wire [35:0] _GEN_30; // @[TensorUtil.scala 277:33:@1394.4]
  wire [35:0] xfer_init_addr; // @[TensorUtil.scala 277:33:@1394.4]
  wire [32:0] _T_162; // @[TensorUtil.scala 278:31:@1395.4]
  wire [31:0] xfer_split_addr; // @[TensorUtil.scala 278:31:@1396.4]
  wire [31:0] _GEN_31; // @[TensorUtil.scala 279:32:@1397.4]
  wire [32:0] _T_163; // @[TensorUtil.scala 279:32:@1397.4]
  wire [31:0] xfer_stride_addr; // @[TensorUtil.scala 279:32:@1398.4]
  wire [35:0] _GEN_12; // @[TensorUtil.scala 281:55:@1399.4]
  wire [11:0] _T_164; // @[TensorUtil.scala 281:55:@1399.4]
  wire [12:0] _T_165; // @[TensorUtil.scala 281:38:@1400.4]
  wire [12:0] _T_166; // @[TensorUtil.scala 281:38:@1401.4]
  wire [11:0] xfer_init_bytes; // @[TensorUtil.scala 281:38:@1402.4]
  wire [8:0] xfer_init_pulses; // @[TensorUtil.scala 282:43:@1403.4]
  wire [31:0] _GEN_16; // @[TensorUtil.scala 283:56:@1404.4]
  wire [11:0] _T_167; // @[TensorUtil.scala 283:56:@1404.4]
  wire [12:0] _T_168; // @[TensorUtil.scala 283:38:@1405.4]
  wire [12:0] _T_169; // @[TensorUtil.scala 283:38:@1406.4]
  wire [11:0] xfer_split_bytes; // @[TensorUtil.scala 283:38:@1407.4]
  wire [8:0] xfer_split_pulses; // @[TensorUtil.scala 284:44:@1408.4]
  wire [31:0] _GEN_18; // @[TensorUtil.scala 285:57:@1409.4]
  wire [11:0] _T_170; // @[TensorUtil.scala 285:57:@1409.4]
  wire [12:0] _T_171; // @[TensorUtil.scala 285:38:@1410.4]
  wire [12:0] _T_172; // @[TensorUtil.scala 285:38:@1411.4]
  wire [11:0] xfer_stride_bytes; // @[TensorUtil.scala 285:38:@1412.4]
  wire [8:0] xfer_stride_pulses; // @[TensorUtil.scala 286:45:@1413.4]
  wire  _T_173; // @[TensorUtil.scala 288:21:@1414.4]
  wire  _T_175; // @[TensorUtil.scala 289:10:@1415.4]
  wire  _T_176; // @[TensorUtil.scala 288:29:@1416.4]
  wire [16:0] _T_178; // @[TensorUtil.scala 290:24:@1417.4]
  wire [16:0] _T_179; // @[TensorUtil.scala 290:24:@1418.4]
  wire [15:0] _T_180; // @[TensorUtil.scala 290:24:@1419.4]
  wire  _T_181; // @[TensorUtil.scala 290:10:@1420.4]
  wire  stride; // @[TensorUtil.scala 289:18:@1421.4]
  wire  _T_184; // @[TensorUtil.scala 292:35:@1423.4]
  wire  split; // @[TensorUtil.scala 292:28:@1424.4]
  wire [16:0] _GEN_32; // @[TensorUtil.scala 296:16:@1427.6]
  wire  _T_185; // @[TensorUtil.scala 296:16:@1427.6]
  wire [9:0] _T_188; // @[TensorUtil.scala 300:31:@1433.8]
  wire [9:0] _T_189; // @[TensorUtil.scala 300:31:@1434.8]
  wire [8:0] _T_190; // @[TensorUtil.scala 300:31:@1435.8]
  wire [17:0] _T_191; // @[TensorUtil.scala 301:21:@1437.8]
  wire [17:0] _T_192; // @[TensorUtil.scala 301:21:@1438.8]
  wire [16:0] _T_193; // @[TensorUtil.scala 301:21:@1439.8]
  wire [16:0] _GEN_0; // @[TensorUtil.scala 296:36:@1428.6]
  wire [16:0] _GEN_1; // @[TensorUtil.scala 296:36:@1428.6]
  wire  _T_194; // @[TensorUtil.scala 303:25:@1444.6]
  wire [16:0] _GEN_34; // @[TensorUtil.scala 305:16:@1447.8]
  wire  _T_195; // @[TensorUtil.scala 305:16:@1447.8]
  wire [9:0] _T_198; // @[TensorUtil.scala 309:33:@1453.10]
  wire [9:0] _T_199; // @[TensorUtil.scala 309:33:@1454.10]
  wire [8:0] _T_200; // @[TensorUtil.scala 309:33:@1455.10]
  wire [17:0] _T_201; // @[TensorUtil.scala 310:21:@1457.10]
  wire [17:0] _T_202; // @[TensorUtil.scala 310:21:@1458.10]
  wire [16:0] _T_203; // @[TensorUtil.scala 310:21:@1459.10]
  wire [16:0] _GEN_2; // @[TensorUtil.scala 305:38:@1448.8]
  wire [16:0] _GEN_3; // @[TensorUtil.scala 305:38:@1448.8]
  wire  _T_204; // @[TensorUtil.scala 312:25:@1464.8]
  wire [15:0] _GEN_36; // @[TensorUtil.scala 314:15:@1467.10]
  wire  _T_205; // @[TensorUtil.scala 314:15:@1467.10]
  wire [9:0] _T_208; // @[TensorUtil.scala 318:32:@1473.12]
  wire [9:0] _T_209; // @[TensorUtil.scala 318:32:@1474.12]
  wire [8:0] _T_210; // @[TensorUtil.scala 318:32:@1475.12]
  wire [16:0] _T_211; // @[TensorUtil.scala 319:20:@1477.12]
  wire [16:0] _T_212; // @[TensorUtil.scala 319:20:@1478.12]
  wire [15:0] _T_213; // @[TensorUtil.scala 319:20:@1479.12]
  wire [15:0] _GEN_4; // @[TensorUtil.scala 314:36:@1468.10]
  wire [15:0] _GEN_5; // @[TensorUtil.scala 314:36:@1468.10]
  wire [31:0] _GEN_6; // @[TensorUtil.scala 312:35:@1465.8]
  wire [15:0] _GEN_7; // @[TensorUtil.scala 312:35:@1465.8]
  wire [15:0] _GEN_8; // @[TensorUtil.scala 312:35:@1465.8]
  wire [31:0] _GEN_9; // @[TensorUtil.scala 303:36:@1445.6]
  wire [16:0] _GEN_10; // @[TensorUtil.scala 303:36:@1445.6]
  wire [16:0] _GEN_11; // @[TensorUtil.scala 303:36:@1445.6]
  wire [16:0] _GEN_13; // @[TensorUtil.scala 294:18:@1425.4]
  wire [16:0] _GEN_14; // @[TensorUtil.scala 294:18:@1425.4]
  wire [8:0] _T_216; // @[TensorUtil.scala 326:18:@1488.8]
  wire [7:0] _T_217; // @[TensorUtil.scala 326:18:@1489.8]
  wire [7:0] _GEN_15; // @[TensorUtil.scala 325:26:@1487.6]
  wire  _T_219; // @[TensorUtil.scala 331:25:@1496.6]
  wire [16:0] _T_221; // @[TensorUtil.scala 332:18:@1498.8]
  wire [15:0] _T_222; // @[TensorUtil.scala 332:18:@1499.8]
  wire [15:0] _GEN_17; // @[TensorUtil.scala 331:36:@1497.6]
  wire [31:0] _GEN_19; // @[TensorUtil.scala 341:24:@1512.10]
  wire [31:0] _GEN_20; // @[TensorUtil.scala 341:24:@1512.10]
  wire [31:0] _GEN_21; // @[TensorUtil.scala 339:17:@1508.8]
  wire [31:0] _GEN_22; // @[TensorUtil.scala 339:17:@1508.8]
  wire [31:0] _GEN_23; // @[TensorUtil.scala 338:26:@1507.6]
  wire [31:0] _GEN_24; // @[TensorUtil.scala 338:26:@1507.6]
  wire [35:0] _GEN_25; // @[TensorUtil.scala 335:18:@1502.4]
  wire [35:0] _GEN_26; // @[TensorUtil.scala 335:18:@1502.4]
  wire  _T_232; // @[TensorUtil.scala 354:10:@1529.4]
  assign dec_dram_offset = io_inst[56:25]; // @[TensorUtil.scala 251:29:@1298.4]
  assign dec_ysize = io_inst[79:64]; // @[TensorUtil.scala 251:29:@1302.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 251:29:@1304.4]
  assign dec_xstride = io_inst[111:96]; // @[TensorUtil.scala 251:29:@1306.4]
  assign _GEN_27 = {{1'd0}, dec_xsize}; // @[TensorUtil.scala 269:26:@1385.4]
  assign _T_154 = _GEN_27 << 1; // @[TensorUtil.scala 269:26:@1385.4]
  assign _T_156 = _T_154 - 17'h1; // @[TensorUtil.scala 269:51:@1386.4]
  assign _T_157 = $unsigned(_T_156); // @[TensorUtil.scala 269:51:@1387.4]
  assign xsize = _T_157[16:0]; // @[TensorUtil.scala 269:51:@1388.4]
  assign _GEN_28 = {{4'd0}, dec_xstride}; // @[TensorUtil.scala 275:35:@1391.4]
  assign xstride_bytes = _GEN_28 << 4; // @[TensorUtil.scala 275:35:@1391.4]
  assign _GEN_29 = {{4'd0}, dec_dram_offset}; // @[TensorUtil.scala 277:66:@1392.4]
  assign _T_160 = _GEN_29 << 4; // @[TensorUtil.scala 277:66:@1392.4]
  assign _T_161 = 36'hffffffff & _T_160; // @[TensorUtil.scala 277:47:@1393.4]
  assign _GEN_30 = {{4'd0}, io_baddr}; // @[TensorUtil.scala 277:33:@1394.4]
  assign xfer_init_addr = _GEN_30 | _T_161; // @[TensorUtil.scala 277:33:@1394.4]
  assign _T_162 = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@1395.4]
  assign xfer_split_addr = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@1396.4]
  assign _GEN_31 = {{12'd0}, xstride_bytes}; // @[TensorUtil.scala 279:32:@1397.4]
  assign _T_163 = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@1397.4]
  assign xfer_stride_addr = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@1398.4]
  assign _GEN_12 = xfer_init_addr % 36'h800; // @[TensorUtil.scala 281:55:@1399.4]
  assign _T_164 = _GEN_12[11:0]; // @[TensorUtil.scala 281:55:@1399.4]
  assign _T_165 = 12'h800 - _T_164; // @[TensorUtil.scala 281:38:@1400.4]
  assign _T_166 = $unsigned(_T_165); // @[TensorUtil.scala 281:38:@1401.4]
  assign xfer_init_bytes = _T_166[11:0]; // @[TensorUtil.scala 281:38:@1402.4]
  assign xfer_init_pulses = xfer_init_bytes[11:3]; // @[TensorUtil.scala 282:43:@1403.4]
  assign _GEN_16 = xfer_split_addr % 32'h800; // @[TensorUtil.scala 283:56:@1404.4]
  assign _T_167 = _GEN_16[11:0]; // @[TensorUtil.scala 283:56:@1404.4]
  assign _T_168 = 12'h800 - _T_167; // @[TensorUtil.scala 283:38:@1405.4]
  assign _T_169 = $unsigned(_T_168); // @[TensorUtil.scala 283:38:@1406.4]
  assign xfer_split_bytes = _T_169[11:0]; // @[TensorUtil.scala 283:38:@1407.4]
  assign xfer_split_pulses = xfer_split_bytes[11:3]; // @[TensorUtil.scala 284:44:@1408.4]
  assign _GEN_18 = xfer_stride_addr % 32'h800; // @[TensorUtil.scala 285:57:@1409.4]
  assign _T_170 = _GEN_18[11:0]; // @[TensorUtil.scala 285:57:@1409.4]
  assign _T_171 = 12'h800 - _T_170; // @[TensorUtil.scala 285:38:@1410.4]
  assign _T_172 = $unsigned(_T_171); // @[TensorUtil.scala 285:38:@1411.4]
  assign xfer_stride_bytes = _T_172[11:0]; // @[TensorUtil.scala 285:38:@1412.4]
  assign xfer_stride_pulses = xfer_stride_bytes[11:3]; // @[TensorUtil.scala 286:45:@1413.4]
  assign _T_173 = xcnt == len; // @[TensorUtil.scala 288:21:@1414.4]
  assign _T_175 = xrem == 16'h0; // @[TensorUtil.scala 289:10:@1415.4]
  assign _T_176 = _T_173 & _T_175; // @[TensorUtil.scala 288:29:@1416.4]
  assign _T_178 = dec_ysize - 16'h1; // @[TensorUtil.scala 290:24:@1417.4]
  assign _T_179 = $unsigned(_T_178); // @[TensorUtil.scala 290:24:@1418.4]
  assign _T_180 = _T_179[15:0]; // @[TensorUtil.scala 290:24:@1419.4]
  assign _T_181 = ycnt != _T_180; // @[TensorUtil.scala 290:10:@1420.4]
  assign stride = _T_176 & _T_181; // @[TensorUtil.scala 289:18:@1421.4]
  assign _T_184 = xrem != 16'h0; // @[TensorUtil.scala 292:35:@1423.4]
  assign split = _T_173 & _T_184; // @[TensorUtil.scala 292:28:@1424.4]
  assign _GEN_32 = {{8'd0}, xfer_init_pulses}; // @[TensorUtil.scala 296:16:@1427.6]
  assign _T_185 = xsize < _GEN_32; // @[TensorUtil.scala 296:16:@1427.6]
  assign _T_188 = xfer_init_pulses - 9'h1; // @[TensorUtil.scala 300:31:@1433.8]
  assign _T_189 = $unsigned(_T_188); // @[TensorUtil.scala 300:31:@1434.8]
  assign _T_190 = _T_189[8:0]; // @[TensorUtil.scala 300:31:@1435.8]
  assign _T_191 = xsize - _GEN_32; // @[TensorUtil.scala 301:21:@1437.8]
  assign _T_192 = $unsigned(_T_191); // @[TensorUtil.scala 301:21:@1438.8]
  assign _T_193 = _T_192[16:0]; // @[TensorUtil.scala 301:21:@1439.8]
  assign _GEN_0 = _T_185 ? xsize : {{8'd0}, _T_190}; // @[TensorUtil.scala 296:36:@1428.6]
  assign _GEN_1 = _T_185 ? 17'h0 : _T_193; // @[TensorUtil.scala 296:36:@1428.6]
  assign _T_194 = io_xupdate & stride; // @[TensorUtil.scala 303:25:@1444.6]
  assign _GEN_34 = {{8'd0}, xfer_stride_pulses}; // @[TensorUtil.scala 305:16:@1447.8]
  assign _T_195 = xsize < _GEN_34; // @[TensorUtil.scala 305:16:@1447.8]
  assign _T_198 = xfer_stride_pulses - 9'h1; // @[TensorUtil.scala 309:33:@1453.10]
  assign _T_199 = $unsigned(_T_198); // @[TensorUtil.scala 309:33:@1454.10]
  assign _T_200 = _T_199[8:0]; // @[TensorUtil.scala 309:33:@1455.10]
  assign _T_201 = xsize - _GEN_34; // @[TensorUtil.scala 310:21:@1457.10]
  assign _T_202 = $unsigned(_T_201); // @[TensorUtil.scala 310:21:@1458.10]
  assign _T_203 = _T_202[16:0]; // @[TensorUtil.scala 310:21:@1459.10]
  assign _GEN_2 = _T_195 ? xsize : {{8'd0}, _T_200}; // @[TensorUtil.scala 305:38:@1448.8]
  assign _GEN_3 = _T_195 ? 17'h0 : _T_203; // @[TensorUtil.scala 305:38:@1448.8]
  assign _T_204 = io_xupdate & split; // @[TensorUtil.scala 312:25:@1464.8]
  assign _GEN_36 = {{7'd0}, xfer_split_pulses}; // @[TensorUtil.scala 314:15:@1467.10]
  assign _T_205 = xrem < _GEN_36; // @[TensorUtil.scala 314:15:@1467.10]
  assign _T_208 = xfer_split_pulses - 9'h1; // @[TensorUtil.scala 318:32:@1473.12]
  assign _T_209 = $unsigned(_T_208); // @[TensorUtil.scala 318:32:@1474.12]
  assign _T_210 = _T_209[8:0]; // @[TensorUtil.scala 318:32:@1475.12]
  assign _T_211 = xrem - _GEN_36; // @[TensorUtil.scala 319:20:@1477.12]
  assign _T_212 = $unsigned(_T_211); // @[TensorUtil.scala 319:20:@1478.12]
  assign _T_213 = _T_212[15:0]; // @[TensorUtil.scala 319:20:@1479.12]
  assign _GEN_4 = _T_205 ? xrem : {{7'd0}, _T_210}; // @[TensorUtil.scala 314:36:@1468.10]
  assign _GEN_5 = _T_205 ? 16'h0 : _T_213; // @[TensorUtil.scala 314:36:@1468.10]
  assign _GEN_6 = _T_204 ? {{20'd0}, xfer_split_bytes} : xfer_bytes; // @[TensorUtil.scala 312:35:@1465.8]
  assign _GEN_7 = _T_204 ? _GEN_4 : {{8'd0}, len}; // @[TensorUtil.scala 312:35:@1465.8]
  assign _GEN_8 = _T_204 ? _GEN_5 : xrem; // @[TensorUtil.scala 312:35:@1465.8]
  assign _GEN_9 = _T_194 ? {{20'd0}, xfer_stride_bytes} : _GEN_6; // @[TensorUtil.scala 303:36:@1445.6]
  assign _GEN_10 = _T_194 ? _GEN_2 : {{1'd0}, _GEN_7}; // @[TensorUtil.scala 303:36:@1445.6]
  assign _GEN_11 = _T_194 ? _GEN_3 : {{1'd0}, _GEN_8}; // @[TensorUtil.scala 303:36:@1445.6]
  assign _GEN_13 = io_start ? _GEN_0 : _GEN_10; // @[TensorUtil.scala 294:18:@1425.4]
  assign _GEN_14 = io_start ? _GEN_1 : _GEN_11; // @[TensorUtil.scala 294:18:@1425.4]
  assign _T_216 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@1488.8]
  assign _T_217 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@1489.8]
  assign _GEN_15 = io_xupdate ? _T_217 : xcnt; // @[TensorUtil.scala 325:26:@1487.6]
  assign _T_219 = io_yupdate & stride; // @[TensorUtil.scala 331:25:@1496.6]
  assign _T_221 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@1498.8]
  assign _T_222 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@1499.8]
  assign _GEN_17 = _T_219 ? _T_222 : ycnt; // @[TensorUtil.scala 331:36:@1497.6]
  assign _GEN_19 = stride ? xfer_stride_addr : caddr; // @[TensorUtil.scala 341:24:@1512.10]
  assign _GEN_20 = stride ? xfer_stride_addr : baddr; // @[TensorUtil.scala 341:24:@1512.10]
  assign _GEN_21 = split ? xfer_split_addr : _GEN_19; // @[TensorUtil.scala 339:17:@1508.8]
  assign _GEN_22 = split ? baddr : _GEN_20; // @[TensorUtil.scala 339:17:@1508.8]
  assign _GEN_23 = io_yupdate ? _GEN_21 : caddr; // @[TensorUtil.scala 338:26:@1507.6]
  assign _GEN_24 = io_yupdate ? _GEN_22 : baddr; // @[TensorUtil.scala 338:26:@1507.6]
  assign _GEN_25 = io_start ? xfer_init_addr : {{4'd0}, _GEN_23}; // @[TensorUtil.scala 335:18:@1502.4]
  assign _GEN_26 = io_start ? xfer_init_addr : {{4'd0}, _GEN_24}; // @[TensorUtil.scala 335:18:@1502.4]
  assign _T_232 = ycnt == _T_180; // @[TensorUtil.scala 354:10:@1529.4]
  assign io_done = _T_176 & _T_232; // @[TensorUtil.scala 352:11:@1531.4]
  assign io_stride = _T_176 & _T_181; // @[TensorUtil.scala 347:13:@1517.4]
  assign io_split = _T_173 & _T_184; // @[TensorUtil.scala 348:12:@1518.4]
  assign io_addr = caddr; // @[TensorUtil.scala 350:11:@1521.4]
  assign io_len = len; // @[TensorUtil.scala 351:10:@1522.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  caddr = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  baddr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  len = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  xcnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xrem = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ycnt = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  xfer_bytes = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    caddr <= _GEN_25[31:0];
    baddr <= _GEN_26[31:0];
    len <= _GEN_13[7:0];
    if (io_xinit) begin
      xcnt <= 8'h0;
    end else begin
      if (io_xupdate) begin
        xcnt <= _T_217;
      end
    end
    xrem <= _GEN_14[15:0];
    if (io_start) begin
      ycnt <= 16'h0;
    end else begin
      if (_T_219) begin
        ycnt <= _T_222;
      end
    end
    if (io_start) begin
      xfer_bytes <= {{20'd0}, xfer_init_bytes};
    end else begin
      if (_T_194) begin
        xfer_bytes <= {{20'd0}, xfer_stride_bytes};
      end else begin
        if (_T_204) begin
          xfer_bytes <= {{20'd0}, xfer_split_bytes};
        end
      end
    end
  end
endmodule
module TensorPadCtrl( // @[:@1533.2]
  input          clock, // @[:@1534.4]
  input          reset, // @[:@1535.4]
  input          io_start, // @[:@1536.4]
  output         io_done, // @[:@1536.4]
  input  [127:0] io_inst // @[:@1536.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@1561.4]
  wire [3:0] dec_ypad_0; // @[TensorUtil.scala 173:29:@1565.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@1569.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@1571.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@1573.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@1574.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@1575.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@1576.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@1577.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@1577.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@1578.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@1579.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@1579.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@1580.4]
  wire [16:0] _GEN_12; // @[TensorUtil.scala 182:46:@1581.4]
  wire [16:0] _T_39; // @[TensorUtil.scala 182:46:@1581.4]
  wire [17:0] _T_41; // @[TensorUtil.scala 182:71:@1582.4]
  wire [17:0] _T_42; // @[TensorUtil.scala 182:71:@1583.4]
  wire [16:0] xval; // @[TensorUtil.scala 182:71:@1584.4]
  wire  _T_44; // @[TensorUtil.scala 190:22:@1585.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 190:42:@1586.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 190:42:@1587.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 190:42:@1588.4]
  wire [3:0] yval; // @[TensorUtil.scala 190:10:@1589.4]
  reg  state; // @[TensorUtil.scala 197:22:@1590.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@1591.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@1593.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@1600.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@1601.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@1602.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@1603.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@1599.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@1592.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@1607.4]
  wire [16:0] _GEN_4; // @[TensorUtil.scala 212:25:@1608.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@1614.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@1621.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@1622.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@1620.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@1626.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@1627.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@1634.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@1636.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@1637.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@1635.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@1642.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@1561.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorUtil.scala 173:29:@1565.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@1569.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@1571.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@1577.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@1577.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@1578.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@1579.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@1579.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@1580.4]
  assign _GEN_12 = {{1'd0}, _T_38}; // @[TensorUtil.scala 182:46:@1581.4]
  assign _T_39 = _GEN_12 << 1; // @[TensorUtil.scala 182:46:@1581.4]
  assign _T_41 = _T_39 - 17'h1; // @[TensorUtil.scala 182:71:@1582.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@1583.4]
  assign xval = _T_42[16:0]; // @[TensorUtil.scala 182:71:@1584.4]
  assign _T_44 = dec_ypad_0 != 4'h0; // @[TensorUtil.scala 190:22:@1585.4]
  assign _T_46 = dec_ypad_0 - 4'h1; // @[TensorUtil.scala 190:42:@1586.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 190:42:@1587.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 190:42:@1588.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 190:10:@1589.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@1591.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@1593.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@1600.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@1601.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@1602.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@1603.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@1599.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@1592.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@1607.4]
  assign _GEN_4 = _T_56 ? xval : {{1'd0}, xmax}; // @[TensorUtil.scala 212:25:@1608.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@1614.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1621.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1622.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@1620.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@1626.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@1627.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@1634.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@1636.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@1637.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@1635.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@1642.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@1645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_1( // @[:@1647.2]
  input          clock, // @[:@1648.4]
  input          reset, // @[:@1649.4]
  input          io_start, // @[:@1650.4]
  output         io_done, // @[:@1650.4]
  input  [127:0] io_inst // @[:@1650.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@1675.4]
  wire [3:0] dec_ypad_1; // @[TensorUtil.scala 173:29:@1681.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@1683.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@1685.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@1687.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@1688.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@1689.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@1690.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@1691.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@1691.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@1692.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@1693.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@1693.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@1694.4]
  wire [16:0] _GEN_12; // @[TensorUtil.scala 182:46:@1695.4]
  wire [16:0] _T_39; // @[TensorUtil.scala 182:46:@1695.4]
  wire [17:0] _T_41; // @[TensorUtil.scala 182:71:@1696.4]
  wire [17:0] _T_42; // @[TensorUtil.scala 182:71:@1697.4]
  wire [16:0] xval; // @[TensorUtil.scala 182:71:@1698.4]
  wire  _T_44; // @[TensorUtil.scala 192:22:@1699.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 192:42:@1700.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 192:42:@1701.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 192:42:@1702.4]
  wire [3:0] yval; // @[TensorUtil.scala 192:10:@1703.4]
  reg  state; // @[TensorUtil.scala 197:22:@1704.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@1705.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@1707.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@1714.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@1715.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@1716.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@1717.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@1713.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@1706.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@1721.4]
  wire [16:0] _GEN_4; // @[TensorUtil.scala 212:25:@1722.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@1728.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@1735.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@1736.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@1734.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@1740.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@1741.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@1748.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@1750.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@1751.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@1749.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@1756.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@1675.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorUtil.scala 173:29:@1681.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@1683.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@1685.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@1691.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@1691.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@1692.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@1693.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@1693.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@1694.4]
  assign _GEN_12 = {{1'd0}, _T_38}; // @[TensorUtil.scala 182:46:@1695.4]
  assign _T_39 = _GEN_12 << 1; // @[TensorUtil.scala 182:46:@1695.4]
  assign _T_41 = _T_39 - 17'h1; // @[TensorUtil.scala 182:71:@1696.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@1697.4]
  assign xval = _T_42[16:0]; // @[TensorUtil.scala 182:71:@1698.4]
  assign _T_44 = dec_ypad_1 != 4'h0; // @[TensorUtil.scala 192:22:@1699.4]
  assign _T_46 = dec_ypad_1 - 4'h1; // @[TensorUtil.scala 192:42:@1700.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 192:42:@1701.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 192:42:@1702.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 192:10:@1703.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@1705.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@1707.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@1714.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@1715.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@1716.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@1717.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@1713.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@1706.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@1721.4]
  assign _GEN_4 = _T_56 ? xval : {{1'd0}, xmax}; // @[TensorUtil.scala 212:25:@1722.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@1728.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1735.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1736.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@1734.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@1740.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@1741.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@1748.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@1750.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@1751.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@1749.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@1756.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@1759.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_2( // @[:@1761.2]
  input          clock, // @[:@1762.4]
  input          reset, // @[:@1763.4]
  input          io_start, // @[:@1764.4]
  output         io_done, // @[:@1764.4]
  input  [127:0] io_inst // @[:@1764.4]
);
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@1797.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@1801.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@1803.4]
  reg [31:0] _RAND_1;
  wire [4:0] _GEN_10; // @[TensorUtil.scala 184:19:@1805.4]
  wire [4:0] _T_35; // @[TensorUtil.scala 184:19:@1805.4]
  wire [5:0] _T_37; // @[TensorUtil.scala 184:44:@1806.4]
  wire [5:0] _T_38; // @[TensorUtil.scala 184:44:@1807.4]
  wire [4:0] xval; // @[TensorUtil.scala 184:44:@1808.4]
  reg  state; // @[TensorUtil.scala 197:22:@1809.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@1810.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@1812.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@1820.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@1822.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@1818.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@1811.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@1826.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@1833.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@1840.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@1841.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@1839.6]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@1797.4]
  assign _GEN_10 = {{1'd0}, dec_xpad_0}; // @[TensorUtil.scala 184:19:@1805.4]
  assign _T_35 = _GEN_10 << 1; // @[TensorUtil.scala 184:19:@1805.4]
  assign _T_37 = _T_35 - 5'h1; // @[TensorUtil.scala 184:44:@1806.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 184:44:@1807.4]
  assign xval = _T_38[4:0]; // @[TensorUtil.scala 184:44:@1808.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@1810.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@1812.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@1820.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@1822.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@1818.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@1811.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@1826.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@1833.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1840.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1841.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@1839.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@1864.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{11'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_3( // @[:@1866.2]
  input          clock, // @[:@1867.4]
  input          reset, // @[:@1868.4]
  input          io_start, // @[:@1869.4]
  output         io_done, // @[:@1869.4]
  input  [127:0] io_inst // @[:@1869.4]
);
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@1904.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@1906.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@1908.4]
  reg [31:0] _RAND_1;
  wire [4:0] _GEN_10; // @[TensorUtil.scala 186:19:@1910.4]
  wire [4:0] _T_35; // @[TensorUtil.scala 186:19:@1910.4]
  wire [5:0] _T_37; // @[TensorUtil.scala 186:44:@1911.4]
  wire [5:0] _T_38; // @[TensorUtil.scala 186:44:@1912.4]
  wire [4:0] xval; // @[TensorUtil.scala 186:44:@1913.4]
  reg  state; // @[TensorUtil.scala 197:22:@1914.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@1915.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@1917.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@1925.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@1927.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@1923.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@1916.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@1931.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@1938.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@1945.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@1946.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@1944.6]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@1904.4]
  assign _GEN_10 = {{1'd0}, dec_xpad_1}; // @[TensorUtil.scala 186:19:@1910.4]
  assign _T_35 = _GEN_10 << 1; // @[TensorUtil.scala 186:19:@1910.4]
  assign _T_37 = _T_35 - 5'h1; // @[TensorUtil.scala 186:44:@1911.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 186:44:@1912.4]
  assign xval = _T_38[4:0]; // @[TensorUtil.scala 186:44:@1913.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@1915.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@1917.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@1925.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@1927.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@1923.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@1916.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@1931.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@1938.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1945.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@1946.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@1944.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@1969.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{11'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorLoad( // @[:@1971.2]
  input          clock, // @[:@1972.4]
  input          reset, // @[:@1973.4]
  input          io_start, // @[:@1974.4]
  output         io_done, // @[:@1974.4]
  input  [127:0] io_inst, // @[:@1974.4]
  input  [31:0]  io_baddr, // @[:@1974.4]
  input          io_vme_rd_cmd_ready, // @[:@1974.4]
  output         io_vme_rd_cmd_valid, // @[:@1974.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@1974.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@1974.4]
  output         io_vme_rd_data_ready, // @[:@1974.4]
  input          io_vme_rd_data_valid, // @[:@1974.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@1974.4]
  input          io_tensor_rd_idx_valid, // @[:@1974.4]
  input  [10:0]  io_tensor_rd_idx_bits, // @[:@1974.4]
  output         io_tensor_rd_data_valid, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_0, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_1, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_2, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_3, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_4, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_5, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_6, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_7, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_8, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_9, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_10, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_11, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_12, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_13, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_14, // @[:@1974.4]
  output [7:0]   io_tensor_rd_data_bits_0_15 // @[:@1974.4]
);
  wire  dataCtrl_clock; // @[TensorLoad.scala 52:24:@2011.4]
  wire  dataCtrl_io_start; // @[TensorLoad.scala 52:24:@2011.4]
  wire  dataCtrl_io_done; // @[TensorLoad.scala 52:24:@2011.4]
  wire [127:0] dataCtrl_io_inst; // @[TensorLoad.scala 52:24:@2011.4]
  wire [31:0] dataCtrl_io_baddr; // @[TensorLoad.scala 52:24:@2011.4]
  wire  dataCtrl_io_xinit; // @[TensorLoad.scala 52:24:@2011.4]
  wire  dataCtrl_io_xupdate; // @[TensorLoad.scala 52:24:@2011.4]
  wire  dataCtrl_io_yupdate; // @[TensorLoad.scala 52:24:@2011.4]
  wire  dataCtrl_io_stride; // @[TensorLoad.scala 52:24:@2011.4]
  wire  dataCtrl_io_split; // @[TensorLoad.scala 52:24:@2011.4]
  wire [31:0] dataCtrl_io_addr; // @[TensorLoad.scala 52:24:@2011.4]
  wire [7:0] dataCtrl_io_len; // @[TensorLoad.scala 52:24:@2011.4]
  wire  yPadCtrl0_clock; // @[TensorLoad.scala 55:25:@2015.4]
  wire  yPadCtrl0_reset; // @[TensorLoad.scala 55:25:@2015.4]
  wire  yPadCtrl0_io_start; // @[TensorLoad.scala 55:25:@2015.4]
  wire  yPadCtrl0_io_done; // @[TensorLoad.scala 55:25:@2015.4]
  wire [127:0] yPadCtrl0_io_inst; // @[TensorLoad.scala 55:25:@2015.4]
  wire  yPadCtrl1_clock; // @[TensorLoad.scala 56:25:@2018.4]
  wire  yPadCtrl1_reset; // @[TensorLoad.scala 56:25:@2018.4]
  wire  yPadCtrl1_io_start; // @[TensorLoad.scala 56:25:@2018.4]
  wire  yPadCtrl1_io_done; // @[TensorLoad.scala 56:25:@2018.4]
  wire [127:0] yPadCtrl1_io_inst; // @[TensorLoad.scala 56:25:@2018.4]
  wire  xPadCtrl0_clock; // @[TensorLoad.scala 57:25:@2021.4]
  wire  xPadCtrl0_reset; // @[TensorLoad.scala 57:25:@2021.4]
  wire  xPadCtrl0_io_start; // @[TensorLoad.scala 57:25:@2021.4]
  wire  xPadCtrl0_io_done; // @[TensorLoad.scala 57:25:@2021.4]
  wire [127:0] xPadCtrl0_io_inst; // @[TensorLoad.scala 57:25:@2021.4]
  wire  xPadCtrl1_clock; // @[TensorLoad.scala 58:25:@2024.4]
  wire  xPadCtrl1_reset; // @[TensorLoad.scala 58:25:@2024.4]
  wire  xPadCtrl1_io_start; // @[TensorLoad.scala 58:25:@2024.4]
  wire  xPadCtrl1_io_done; // @[TensorLoad.scala 58:25:@2024.4]
  wire [127:0] xPadCtrl1_io_inst; // @[TensorLoad.scala 58:25:@2024.4]
  reg [63:0] tensorFile_0_0 [0:2047]; // @[TensorLoad.scala 222:16:@2294.4]
  reg [63:0] _RAND_0;
  wire [63:0] tensorFile_0_0_rdata_0_data; // @[TensorLoad.scala 222:16:@2294.4]
  wire [10:0] tensorFile_0_0_rdata_0_addr; // @[TensorLoad.scala 222:16:@2294.4]
  wire [63:0] tensorFile_0_0__T_866_data; // @[TensorLoad.scala 222:16:@2294.4]
  wire [10:0] tensorFile_0_0__T_866_addr; // @[TensorLoad.scala 222:16:@2294.4]
  wire  tensorFile_0_0__T_866_mask; // @[TensorLoad.scala 222:16:@2294.4]
  wire  tensorFile_0_0__T_866_en; // @[TensorLoad.scala 222:16:@2294.4]
  reg [63:0] tensorFile_0_1 [0:2047]; // @[TensorLoad.scala 222:16:@2294.4]
  reg [63:0] _RAND_1;
  wire [63:0] tensorFile_0_1_rdata_0_data; // @[TensorLoad.scala 222:16:@2294.4]
  wire [10:0] tensorFile_0_1_rdata_0_addr; // @[TensorLoad.scala 222:16:@2294.4]
  wire [63:0] tensorFile_0_1__T_866_data; // @[TensorLoad.scala 222:16:@2294.4]
  wire [10:0] tensorFile_0_1__T_866_addr; // @[TensorLoad.scala 222:16:@2294.4]
  wire  tensorFile_0_1__T_866_mask; // @[TensorLoad.scala 222:16:@2294.4]
  wire  tensorFile_0_1__T_866_en; // @[TensorLoad.scala 222:16:@2294.4]
  wire [15:0] dec_sram_offset; // @[TensorLoad.scala 51:29:@1991.4]
  wire [15:0] dec_xsize; // @[TensorLoad.scala 51:29:@1999.4]
  wire [3:0] dec_ypad_0; // @[TensorLoad.scala 51:29:@2003.4]
  wire [3:0] dec_ypad_1; // @[TensorLoad.scala 51:29:@2005.4]
  wire [3:0] dec_xpad_0; // @[TensorLoad.scala 51:29:@2007.4]
  wire [3:0] dec_xpad_1; // @[TensorLoad.scala 51:29:@2009.4]
  reg  dataCtrlDone; // @[TensorLoad.scala 54:29:@2014.4]
  reg [31:0] _RAND_2;
  reg  tag; // @[TensorLoad.scala 60:16:@2027.4]
  reg [31:0] _RAND_3;
  reg [2:0] state; // @[TensorLoad.scala 65:22:@2029.4]
  reg [31:0] _RAND_4;
  wire  _T_614; // @[Conditional.scala 37:30:@2030.4]
  wire  _T_616; // @[TensorLoad.scala 71:25:@2033.8]
  wire  _T_618; // @[TensorLoad.scala 73:31:@2038.10]
  wire [2:0] _GEN_0; // @[TensorLoad.scala 73:40:@2039.10]
  wire [2:0] _GEN_1; // @[TensorLoad.scala 71:34:@2034.8]
  wire [2:0] _GEN_2; // @[TensorLoad.scala 70:22:@2032.6]
  wire  _T_619; // @[Conditional.scala 37:30:@2048.6]
  wire [2:0] _GEN_4; // @[TensorLoad.scala 81:31:@2050.8]
  wire  _T_622; // @[Conditional.scala 37:30:@2061.8]
  wire [2:0] _GEN_5; // @[TensorLoad.scala 90:31:@2063.10]
  wire  _T_623; // @[Conditional.scala 37:30:@2068.10]
  wire [2:0] _GEN_6; // @[TensorLoad.scala 95:33:@2070.12]
  wire  _T_624; // @[Conditional.scala 37:30:@2075.12]
  wire  _T_626; // @[TensorLoad.scala 102:27:@2079.18]
  wire  _T_628; // @[TensorLoad.scala 104:33:@2084.20]
  wire [2:0] _GEN_7; // @[TensorLoad.scala 104:42:@2085.20]
  wire [2:0] _GEN_8; // @[TensorLoad.scala 102:36:@2080.18]
  wire [2:0] _GEN_10; // @[TensorLoad.scala 110:36:@2095.20]
  wire [2:0] _GEN_11; // @[TensorLoad.scala 117:39:@2108.20]
  wire [2:0] _GEN_12; // @[TensorLoad.scala 109:40:@2093.18]
  wire [2:0] _GEN_13; // @[TensorLoad.scala 101:32:@2078.16]
  wire [2:0] _GEN_14; // @[TensorLoad.scala 100:34:@2077.14]
  wire  _T_633; // @[Conditional.scala 37:30:@2114.14]
  wire [2:0] _GEN_17; // @[TensorLoad.scala 124:28:@2117.18]
  wire [2:0] _GEN_18; // @[TensorLoad.scala 123:31:@2116.16]
  wire  _T_638; // @[Conditional.scala 37:30:@2138.16]
  wire  _T_639; // @[TensorLoad.scala 140:30:@2140.18]
  wire [2:0] _GEN_19; // @[TensorLoad.scala 140:47:@2141.18]
  wire [2:0] _GEN_20; // @[Conditional.scala 39:67:@2139.16]
  wire [2:0] _GEN_21; // @[Conditional.scala 39:67:@2115.14]
  wire [2:0] _GEN_22; // @[Conditional.scala 39:67:@2076.12]
  wire [2:0] _GEN_23; // @[Conditional.scala 39:67:@2069.10]
  wire [2:0] _GEN_24; // @[Conditional.scala 39:67:@2062.8]
  wire [2:0] _GEN_25; // @[Conditional.scala 39:67:@2049.6]
  wire [2:0] _GEN_26; // @[Conditional.scala 40:58:@2031.4]
  wire  _T_640; // @[TensorLoad.scala 147:30:@2145.4]
  wire  _T_641; // @[TensorLoad.scala 147:40:@2146.4]
  wire  _T_643; // @[Decoupled.scala 37:37:@2152.4]
  wire  _T_648; // @[TensorLoad.scala 156:36:@2162.6]
  wire  _GEN_27; // @[TensorLoad.scala 156:57:@2163.6]
  wire  _GEN_28; // @[TensorLoad.scala 154:25:@2157.4]
  wire  _T_653; // @[TensorLoad.scala 161:44:@2168.4]
  wire  _T_660; // @[TensorLoad.scala 164:61:@2174.4]
  wire  _T_661; // @[TensorLoad.scala 164:48:@2175.4]
  wire  _T_662; // @[TensorLoad.scala 165:14:@2176.4]
  wire  _T_663; // @[TensorLoad.scala 165:25:@2177.4]
  wire  _T_664; // @[TensorLoad.scala 165:45:@2178.4]
  wire  _T_665; // @[TensorLoad.scala 164:70:@2179.4]
  wire  _T_671; // @[TensorLoad.scala 169:14:@2185.4]
  wire  _T_672; // @[TensorLoad.scala 169:25:@2186.4]
  wire  _T_673; // @[TensorLoad.scala 168:35:@2187.4]
  wire  _T_675; // @[TensorLoad.scala 170:32:@2189.4]
  wire  _T_676; // @[TensorLoad.scala 170:30:@2190.4]
  wire  _T_677; // @[TensorLoad.scala 170:46:@2191.4]
  wire  _T_680; // @[TensorLoad.scala 170:67:@2193.4]
  wire  _T_681; // @[TensorLoad.scala 169:46:@2194.4]
  wire  _T_685; // @[TensorLoad.scala 171:45:@2198.4]
  wire  _T_686; // @[TensorLoad.scala 170:89:@2199.4]
  wire  _T_691; // @[TensorLoad.scala 173:44:@2204.4]
  wire  _T_692; // @[TensorLoad.scala 174:28:@2205.4]
  wire  _T_693; // @[TensorLoad.scala 174:46:@2206.4]
  wire  _T_696; // @[TensorLoad.scala 174:67:@2208.4]
  wire  _T_697; // @[TensorLoad.scala 174:25:@2209.4]
  wire  _T_699; // @[TensorLoad.scala 182:32:@2216.4]
  wire  _T_702; // @[TensorLoad.scala 190:11:@2223.4]
  wire  _T_703; // @[TensorLoad.scala 189:36:@2224.4]
  wire  _T_705; // @[TensorLoad.scala 190:22:@2226.4]
  wire  _T_706; // @[TensorLoad.scala 192:11:@2227.4]
  wire  isZeroPad; // @[TensorLoad.scala 191:22:@2228.4]
  wire  _T_709; // @[TensorLoad.scala 194:24:@2231.4]
  wire  _T_712; // @[TensorLoad.scala 194:46:@2233.4]
  wire  _T_715; // @[TensorLoad.scala 196:36:@2239.6]
  wire [1:0] _T_717; // @[TensorLoad.scala 197:16:@2241.8]
  wire  _T_718; // @[TensorLoad.scala 197:16:@2242.8]
  wire  _GEN_29; // @[TensorLoad.scala 196:50:@2240.6]
  wire  _T_732; // @[TensorLoad.scala 202:51:@2258.6]
  reg [10:0] waddr_cur; // @[TensorLoad.scala 206:22:@2264.4]
  reg [31:0] _RAND_5;
  reg [10:0] waddr_nxt; // @[TensorLoad.scala 207:22:@2265.4]
  reg [31:0] _RAND_6;
  wire [11:0] _T_748; // @[TensorLoad.scala 215:28:@2279.8]
  wire [10:0] _T_749; // @[TensorLoad.scala 215:28:@2280.8]
  wire  _T_751; // @[TensorLoad.scala 216:33:@2285.8]
  wire [15:0] _GEN_66; // @[TensorLoad.scala 217:28:@2287.10]
  wire [16:0] _T_752; // @[TensorLoad.scala 217:28:@2287.10]
  wire [15:0] _T_753; // @[TensorLoad.scala 217:28:@2288.10]
  wire [15:0] _GEN_33; // @[TensorLoad.scala 216:59:@2286.8]
  wire [15:0] _GEN_34; // @[TensorLoad.scala 216:59:@2286.8]
  wire [15:0] _GEN_35; // @[TensorLoad.scala 214:3:@2278.6]
  wire [15:0] _GEN_36; // @[TensorLoad.scala 214:3:@2278.6]
  wire [15:0] _GEN_37; // @[TensorLoad.scala 208:25:@2267.4]
  wire [15:0] _GEN_38; // @[TensorLoad.scala 208:25:@2267.4]
  wire  wmask_0_0; // @[TensorLoad.scala 235:26:@2300.4]
  wire [63:0] wdata_0_0; // @[TensorLoad.scala 236:25:@2302.4]
  reg  rvalid; // @[TensorLoad.scala 252:23:@2351.4]
  reg [31:0] _RAND_7;
  wire  _GEN_51; // @[TensorLoad.scala 256:26:@2356.4]
  wire [127:0] _T_887; // @[TensorLoad.scala 259:38:@2362.4]
  wire  _T_1035; // @[TensorLoad.scala 263:96:@2418.4]
  wire  done_no_pad; // @[TensorLoad.scala 263:83:@2419.4]
  wire  done_x_pad; // @[TensorLoad.scala 264:72:@2424.4]
  wire  _T_1042; // @[TensorLoad.scala 265:37:@2426.4]
  wire  done_y_pad; // @[TensorLoad.scala 265:52:@2427.4]
  wire  _T_1043; // @[TensorLoad.scala 266:26:@2428.4]
  reg [10:0] tensorFile_0_0_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [10:0] tensorFile_0_1_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_9;
  TensorDataCtrl dataCtrl ( // @[TensorLoad.scala 52:24:@2011.4]
    .clock(dataCtrl_clock),
    .io_start(dataCtrl_io_start),
    .io_done(dataCtrl_io_done),
    .io_inst(dataCtrl_io_inst),
    .io_baddr(dataCtrl_io_baddr),
    .io_xinit(dataCtrl_io_xinit),
    .io_xupdate(dataCtrl_io_xupdate),
    .io_yupdate(dataCtrl_io_yupdate),
    .io_stride(dataCtrl_io_stride),
    .io_split(dataCtrl_io_split),
    .io_addr(dataCtrl_io_addr),
    .io_len(dataCtrl_io_len)
  );
  TensorPadCtrl yPadCtrl0 ( // @[TensorLoad.scala 55:25:@2015.4]
    .clock(yPadCtrl0_clock),
    .reset(yPadCtrl0_reset),
    .io_start(yPadCtrl0_io_start),
    .io_done(yPadCtrl0_io_done),
    .io_inst(yPadCtrl0_io_inst)
  );
  TensorPadCtrl_1 yPadCtrl1 ( // @[TensorLoad.scala 56:25:@2018.4]
    .clock(yPadCtrl1_clock),
    .reset(yPadCtrl1_reset),
    .io_start(yPadCtrl1_io_start),
    .io_done(yPadCtrl1_io_done),
    .io_inst(yPadCtrl1_io_inst)
  );
  TensorPadCtrl_2 xPadCtrl0 ( // @[TensorLoad.scala 57:25:@2021.4]
    .clock(xPadCtrl0_clock),
    .reset(xPadCtrl0_reset),
    .io_start(xPadCtrl0_io_start),
    .io_done(xPadCtrl0_io_done),
    .io_inst(xPadCtrl0_io_inst)
  );
  TensorPadCtrl_3 xPadCtrl1 ( // @[TensorLoad.scala 58:25:@2024.4]
    .clock(xPadCtrl1_clock),
    .reset(xPadCtrl1_reset),
    .io_start(xPadCtrl1_io_start),
    .io_done(xPadCtrl1_io_done),
    .io_inst(xPadCtrl1_io_inst)
  );
  assign tensorFile_0_0_rdata_0_addr = tensorFile_0_0_rdata_0_addr_pipe_0;
  assign tensorFile_0_0_rdata_0_data = tensorFile_0_0[tensorFile_0_0_rdata_0_addr]; // @[TensorLoad.scala 222:16:@2294.4]
  assign tensorFile_0_0__T_866_data = _T_640 ? 64'h0 : wdata_0_0;
  assign tensorFile_0_0__T_866_addr = _T_640 ? 11'h0 : waddr_cur;
  assign tensorFile_0_0__T_866_mask = _T_640 ? 1'h1 : wmask_0_0;
  assign tensorFile_0_0__T_866_en = _T_640 ? 1'h0 : _T_715;
  assign tensorFile_0_1_rdata_0_addr = tensorFile_0_1_rdata_0_addr_pipe_0;
  assign tensorFile_0_1_rdata_0_data = tensorFile_0_1[tensorFile_0_1_rdata_0_addr]; // @[TensorLoad.scala 222:16:@2294.4]
  assign tensorFile_0_1__T_866_data = _T_640 ? 64'h0 : wdata_0_0;
  assign tensorFile_0_1__T_866_addr = _T_640 ? 11'h0 : waddr_cur;
  assign tensorFile_0_1__T_866_mask = _T_640 ? 1'h1 : tag;
  assign tensorFile_0_1__T_866_en = _T_640 ? 1'h0 : _T_715;
  assign dec_sram_offset = io_inst[24:9]; // @[TensorLoad.scala 51:29:@1991.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorLoad.scala 51:29:@1999.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorLoad.scala 51:29:@2003.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorLoad.scala 51:29:@2005.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorLoad.scala 51:29:@2007.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorLoad.scala 51:29:@2009.4]
  assign _T_614 = 3'h0 == state; // @[Conditional.scala 37:30:@2030.4]
  assign _T_616 = dec_ypad_0 != 4'h0; // @[TensorLoad.scala 71:25:@2033.8]
  assign _T_618 = dec_xpad_0 != 4'h0; // @[TensorLoad.scala 73:31:@2038.10]
  assign _GEN_0 = _T_618 ? 3'h2 : 3'h3; // @[TensorLoad.scala 73:40:@2039.10]
  assign _GEN_1 = _T_616 ? 3'h1 : _GEN_0; // @[TensorLoad.scala 71:34:@2034.8]
  assign _GEN_2 = io_start ? _GEN_1 : state; // @[TensorLoad.scala 70:22:@2032.6]
  assign _T_619 = 3'h1 == state; // @[Conditional.scala 37:30:@2048.6]
  assign _GEN_4 = yPadCtrl0_io_done ? _GEN_0 : state; // @[TensorLoad.scala 81:31:@2050.8]
  assign _T_622 = 3'h2 == state; // @[Conditional.scala 37:30:@2061.8]
  assign _GEN_5 = xPadCtrl0_io_done ? 3'h3 : state; // @[TensorLoad.scala 90:31:@2063.10]
  assign _T_623 = 3'h3 == state; // @[Conditional.scala 37:30:@2068.10]
  assign _GEN_6 = io_vme_rd_cmd_ready ? 3'h4 : state; // @[TensorLoad.scala 95:33:@2070.12]
  assign _T_624 = 3'h4 == state; // @[Conditional.scala 37:30:@2075.12]
  assign _T_626 = dec_xpad_1 != 4'h0; // @[TensorLoad.scala 102:27:@2079.18]
  assign _T_628 = dec_ypad_1 != 4'h0; // @[TensorLoad.scala 104:33:@2084.20]
  assign _GEN_7 = _T_628 ? 3'h6 : 3'h0; // @[TensorLoad.scala 104:42:@2085.20]
  assign _GEN_8 = _T_626 ? 3'h5 : _GEN_7; // @[TensorLoad.scala 102:36:@2080.18]
  assign _GEN_10 = _T_626 ? 3'h5 : _GEN_0; // @[TensorLoad.scala 110:36:@2095.20]
  assign _GEN_11 = dataCtrl_io_split ? 3'h3 : state; // @[TensorLoad.scala 117:39:@2108.20]
  assign _GEN_12 = dataCtrl_io_stride ? _GEN_10 : _GEN_11; // @[TensorLoad.scala 109:40:@2093.18]
  assign _GEN_13 = dataCtrl_io_done ? _GEN_8 : _GEN_12; // @[TensorLoad.scala 101:32:@2078.16]
  assign _GEN_14 = io_vme_rd_data_valid ? _GEN_13 : state; // @[TensorLoad.scala 100:34:@2077.14]
  assign _T_633 = 3'h5 == state; // @[Conditional.scala 37:30:@2114.14]
  assign _GEN_17 = dataCtrlDone ? _GEN_7 : _GEN_0; // @[TensorLoad.scala 124:28:@2117.18]
  assign _GEN_18 = xPadCtrl1_io_done ? _GEN_17 : state; // @[TensorLoad.scala 123:31:@2116.16]
  assign _T_638 = 3'h6 == state; // @[Conditional.scala 37:30:@2138.16]
  assign _T_639 = yPadCtrl1_io_done & dataCtrlDone; // @[TensorLoad.scala 140:30:@2140.18]
  assign _GEN_19 = _T_639 ? 3'h0 : state; // @[TensorLoad.scala 140:47:@2141.18]
  assign _GEN_20 = _T_638 ? _GEN_19 : state; // @[Conditional.scala 39:67:@2139.16]
  assign _GEN_21 = _T_633 ? _GEN_18 : _GEN_20; // @[Conditional.scala 39:67:@2115.14]
  assign _GEN_22 = _T_624 ? _GEN_14 : _GEN_21; // @[Conditional.scala 39:67:@2076.12]
  assign _GEN_23 = _T_623 ? _GEN_6 : _GEN_22; // @[Conditional.scala 39:67:@2069.10]
  assign _GEN_24 = _T_622 ? _GEN_5 : _GEN_23; // @[Conditional.scala 39:67:@2062.8]
  assign _GEN_25 = _T_619 ? _GEN_4 : _GEN_24; // @[Conditional.scala 39:67:@2049.6]
  assign _GEN_26 = _T_614 ? _GEN_2 : _GEN_25; // @[Conditional.scala 40:58:@2031.4]
  assign _T_640 = state == 3'h0; // @[TensorLoad.scala 147:30:@2145.4]
  assign _T_641 = _T_640 & io_start; // @[TensorLoad.scala 147:40:@2146.4]
  assign _T_643 = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[Decoupled.scala 37:37:@2152.4]
  assign _T_648 = _T_643 & dataCtrl_io_done; // @[TensorLoad.scala 156:36:@2162.6]
  assign _GEN_27 = _T_648 ? 1'h1 : dataCtrlDone; // @[TensorLoad.scala 156:57:@2163.6]
  assign _GEN_28 = _T_640 ? 1'h0 : _GEN_27; // @[TensorLoad.scala 154:25:@2157.4]
  assign _T_653 = _T_616 & _T_640; // @[TensorLoad.scala 161:44:@2168.4]
  assign _T_660 = dec_xpad_1 == 4'h0; // @[TensorLoad.scala 164:61:@2174.4]
  assign _T_661 = _T_648 & _T_660; // @[TensorLoad.scala 164:48:@2175.4]
  assign _T_662 = state == 3'h5; // @[TensorLoad.scala 165:14:@2176.4]
  assign _T_663 = _T_662 & xPadCtrl1_io_done; // @[TensorLoad.scala 165:25:@2177.4]
  assign _T_664 = _T_663 & dataCtrlDone; // @[TensorLoad.scala 165:45:@2178.4]
  assign _T_665 = _T_661 | _T_664; // @[TensorLoad.scala 164:70:@2179.4]
  assign _T_671 = state == 3'h1; // @[TensorLoad.scala 169:14:@2185.4]
  assign _T_672 = _T_671 & yPadCtrl0_io_done; // @[TensorLoad.scala 169:25:@2186.4]
  assign _T_673 = _T_641 | _T_672; // @[TensorLoad.scala 168:35:@2187.4]
  assign _T_675 = ~ dataCtrlDone; // @[TensorLoad.scala 170:32:@2189.4]
  assign _T_676 = _T_643 & _T_675; // @[TensorLoad.scala 170:30:@2190.4]
  assign _T_677 = _T_676 & dataCtrl_io_stride; // @[TensorLoad.scala 170:46:@2191.4]
  assign _T_680 = _T_677 & _T_660; // @[TensorLoad.scala 170:67:@2193.4]
  assign _T_681 = _T_673 | _T_680; // @[TensorLoad.scala 169:46:@2194.4]
  assign _T_685 = _T_663 & _T_675; // @[TensorLoad.scala 171:45:@2198.4]
  assign _T_686 = _T_681 | _T_685; // @[TensorLoad.scala 170:89:@2199.4]
  assign _T_691 = _T_626 & _T_643; // @[TensorLoad.scala 173:44:@2204.4]
  assign _T_692 = ~ dataCtrl_io_done; // @[TensorLoad.scala 174:28:@2205.4]
  assign _T_693 = _T_692 & dataCtrl_io_stride; // @[TensorLoad.scala 174:46:@2206.4]
  assign _T_696 = _T_693 & _T_626; // @[TensorLoad.scala 174:67:@2208.4]
  assign _T_697 = dataCtrl_io_done | _T_696; // @[TensorLoad.scala 174:25:@2209.4]
  assign _T_699 = state == 3'h3; // @[TensorLoad.scala 182:32:@2216.4]
  assign _T_702 = state == 3'h2; // @[TensorLoad.scala 190:11:@2223.4]
  assign _T_703 = _T_671 | _T_702; // @[TensorLoad.scala 189:36:@2224.4]
  assign _T_705 = _T_703 | _T_662; // @[TensorLoad.scala 190:22:@2226.4]
  assign _T_706 = state == 3'h6; // @[TensorLoad.scala 192:11:@2227.4]
  assign isZeroPad = _T_705 | _T_706; // @[TensorLoad.scala 191:22:@2228.4]
  assign _T_709 = _T_640 | _T_699; // @[TensorLoad.scala 194:24:@2231.4]
  assign _T_712 = _T_709 | tag; // @[TensorLoad.scala 194:46:@2233.4]
  assign _T_715 = _T_643 | isZeroPad; // @[TensorLoad.scala 196:36:@2239.6]
  assign _T_717 = tag + 1'h1; // @[TensorLoad.scala 197:16:@2241.8]
  assign _T_718 = tag + 1'h1; // @[TensorLoad.scala 197:16:@2242.8]
  assign _GEN_29 = _T_715 ? _T_718 : tag; // @[TensorLoad.scala 196:50:@2240.6]
  assign _T_732 = _T_715 & tag; // @[TensorLoad.scala 202:51:@2258.6]
  assign _T_748 = waddr_cur + 11'h1; // @[TensorLoad.scala 215:28:@2279.8]
  assign _T_749 = waddr_cur + 11'h1; // @[TensorLoad.scala 215:28:@2280.8]
  assign _T_751 = dataCtrl_io_stride & _T_643; // @[TensorLoad.scala 216:33:@2285.8]
  assign _GEN_66 = {{5'd0}, waddr_nxt}; // @[TensorLoad.scala 217:28:@2287.10]
  assign _T_752 = _GEN_66 + dec_xsize; // @[TensorLoad.scala 217:28:@2287.10]
  assign _T_753 = _GEN_66 + dec_xsize; // @[TensorLoad.scala 217:28:@2288.10]
  assign _GEN_33 = _T_751 ? _T_753 : {{5'd0}, waddr_cur}; // @[TensorLoad.scala 216:59:@2286.8]
  assign _GEN_34 = _T_751 ? _T_753 : {{5'd0}, waddr_nxt}; // @[TensorLoad.scala 216:59:@2286.8]
  assign _GEN_35 = _T_732 ? {{5'd0}, _T_749} : _GEN_33; // @[TensorLoad.scala 214:3:@2278.6]
  assign _GEN_36 = _T_732 ? {{5'd0}, waddr_nxt} : _GEN_34; // @[TensorLoad.scala 214:3:@2278.6]
  assign _GEN_37 = _T_640 ? dec_sram_offset : _GEN_35; // @[TensorLoad.scala 208:25:@2267.4]
  assign _GEN_38 = _T_640 ? dec_sram_offset : _GEN_36; // @[TensorLoad.scala 208:25:@2267.4]
  assign wmask_0_0 = tag == 1'h0; // @[TensorLoad.scala 235:26:@2300.4]
  assign wdata_0_0 = isZeroPad ? 64'h0 : io_vme_rd_data_bits; // @[TensorLoad.scala 236:25:@2302.4]
  assign _GEN_51 = io_tensor_rd_idx_valid; // @[TensorLoad.scala 256:26:@2356.4]
  assign _T_887 = {tensorFile_0_1_rdata_0_data,tensorFile_0_0_rdata_0_data}; // @[TensorLoad.scala 259:38:@2362.4]
  assign _T_1035 = dec_ypad_1 == 4'h0; // @[TensorLoad.scala 263:96:@2418.4]
  assign done_no_pad = _T_661 & _T_1035; // @[TensorLoad.scala 263:83:@2419.4]
  assign done_x_pad = _T_664 & _T_1035; // @[TensorLoad.scala 264:72:@2424.4]
  assign _T_1042 = _T_706 & dataCtrlDone; // @[TensorLoad.scala 265:37:@2426.4]
  assign done_y_pad = _T_1042 & yPadCtrl1_io_done; // @[TensorLoad.scala 265:52:@2427.4]
  assign _T_1043 = done_no_pad | done_x_pad; // @[TensorLoad.scala 266:26:@2428.4]
  assign io_done = _T_1043 | done_y_pad; // @[TensorLoad.scala 266:11:@2430.4]
  assign io_vme_rd_cmd_valid = state == 3'h3; // @[TensorLoad.scala 182:23:@2217.4]
  assign io_vme_rd_cmd_bits_addr = dataCtrl_io_addr; // @[TensorLoad.scala 183:27:@2218.4]
  assign io_vme_rd_cmd_bits_len = dataCtrl_io_len; // @[TensorLoad.scala 184:26:@2219.4]
  assign io_vme_rd_data_ready = state == 3'h4; // @[TensorLoad.scala 186:24:@2221.4]
  assign io_tensor_rd_data_valid = rvalid; // @[TensorLoad.scala 253:27:@2353.4]
  assign io_tensor_rd_data_bits_0_0 = _T_887[7:0]; // @[TensorLoad.scala 259:33:@2398.4]
  assign io_tensor_rd_data_bits_0_1 = _T_887[15:8]; // @[TensorLoad.scala 259:33:@2399.4]
  assign io_tensor_rd_data_bits_0_2 = _T_887[23:16]; // @[TensorLoad.scala 259:33:@2400.4]
  assign io_tensor_rd_data_bits_0_3 = _T_887[31:24]; // @[TensorLoad.scala 259:33:@2401.4]
  assign io_tensor_rd_data_bits_0_4 = _T_887[39:32]; // @[TensorLoad.scala 259:33:@2402.4]
  assign io_tensor_rd_data_bits_0_5 = _T_887[47:40]; // @[TensorLoad.scala 259:33:@2403.4]
  assign io_tensor_rd_data_bits_0_6 = _T_887[55:48]; // @[TensorLoad.scala 259:33:@2404.4]
  assign io_tensor_rd_data_bits_0_7 = _T_887[63:56]; // @[TensorLoad.scala 259:33:@2405.4]
  assign io_tensor_rd_data_bits_0_8 = _T_887[71:64]; // @[TensorLoad.scala 259:33:@2406.4]
  assign io_tensor_rd_data_bits_0_9 = _T_887[79:72]; // @[TensorLoad.scala 259:33:@2407.4]
  assign io_tensor_rd_data_bits_0_10 = _T_887[87:80]; // @[TensorLoad.scala 259:33:@2408.4]
  assign io_tensor_rd_data_bits_0_11 = _T_887[95:88]; // @[TensorLoad.scala 259:33:@2409.4]
  assign io_tensor_rd_data_bits_0_12 = _T_887[103:96]; // @[TensorLoad.scala 259:33:@2410.4]
  assign io_tensor_rd_data_bits_0_13 = _T_887[111:104]; // @[TensorLoad.scala 259:33:@2411.4]
  assign io_tensor_rd_data_bits_0_14 = _T_887[119:112]; // @[TensorLoad.scala 259:33:@2412.4]
  assign io_tensor_rd_data_bits_0_15 = _T_887[127:120]; // @[TensorLoad.scala 259:33:@2413.4]
  assign dataCtrl_clock = clock; // @[:@2012.4]
  assign dataCtrl_io_start = _T_640 & io_start; // @[TensorLoad.scala 147:21:@2147.4]
  assign dataCtrl_io_inst = io_inst; // @[TensorLoad.scala 148:20:@2148.4]
  assign dataCtrl_io_baddr = io_baddr; // @[TensorLoad.scala 149:21:@2149.4]
  assign dataCtrl_io_xinit = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[TensorLoad.scala 150:21:@2151.4]
  assign dataCtrl_io_xupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 151:23:@2153.4]
  assign dataCtrl_io_yupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 152:23:@2155.4]
  assign yPadCtrl0_clock = clock; // @[:@2016.4]
  assign yPadCtrl0_reset = reset; // @[:@2017.4]
  assign yPadCtrl0_io_start = _T_653 & io_start; // @[TensorLoad.scala 161:22:@2170.4]
  assign yPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 176:21:@2212.4]
  assign yPadCtrl1_clock = clock; // @[:@2019.4]
  assign yPadCtrl1_reset = reset; // @[:@2020.4]
  assign yPadCtrl1_io_start = _T_628 & _T_665; // @[TensorLoad.scala 163:22:@2181.4]
  assign yPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 177:21:@2213.4]
  assign xPadCtrl0_clock = clock; // @[:@2022.4]
  assign xPadCtrl0_reset = reset; // @[:@2023.4]
  assign xPadCtrl0_io_start = _T_618 & _T_686; // @[TensorLoad.scala 167:22:@2201.4]
  assign xPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 178:21:@2214.4]
  assign xPadCtrl1_clock = clock; // @[:@2025.4]
  assign xPadCtrl1_reset = reset; // @[:@2026.4]
  assign xPadCtrl1_io_start = _T_691 & _T_697; // @[TensorLoad.scala 173:22:@2211.4]
  assign xPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 179:21:@2215.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_0[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_1[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  dataCtrlDone = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  tag = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  waddr_cur = _RAND_5[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  waddr_nxt = _RAND_6[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rvalid = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tensorFile_0_0_rdata_0_addr_pipe_0 = _RAND_8[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  tensorFile_0_1_rdata_0_addr_pipe_0 = _RAND_9[10:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tensorFile_0_0__T_866_en & tensorFile_0_0__T_866_mask) begin
      tensorFile_0_0[tensorFile_0_0__T_866_addr] <= tensorFile_0_0__T_866_data; // @[TensorLoad.scala 222:16:@2294.4]
    end
    if(tensorFile_0_1__T_866_en & tensorFile_0_1__T_866_mask) begin
      tensorFile_0_1[tensorFile_0_1__T_866_addr] <= tensorFile_0_1__T_866_data; // @[TensorLoad.scala 222:16:@2294.4]
    end
    if (reset) begin
      dataCtrlDone <= 1'h0;
    end else begin
      if (_T_640) begin
        dataCtrlDone <= 1'h0;
      end else begin
        if (_T_648) begin
          dataCtrlDone <= 1'h1;
        end
      end
    end
    if (_T_712) begin
      tag <= 1'h0;
    end else begin
      if (_T_715) begin
        tag <= _T_718;
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_614) begin
        if (io_start) begin
          if (_T_616) begin
            state <= 3'h1;
          end else begin
            if (_T_618) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end
      end else begin
        if (_T_619) begin
          if (yPadCtrl0_io_done) begin
            if (_T_618) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end else begin
          if (_T_622) begin
            if (xPadCtrl0_io_done) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_623) begin
              if (io_vme_rd_cmd_ready) begin
                state <= 3'h4;
              end
            end else begin
              if (_T_624) begin
                if (io_vme_rd_data_valid) begin
                  if (dataCtrl_io_done) begin
                    if (_T_626) begin
                      state <= 3'h5;
                    end else begin
                      if (_T_628) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end
                  end else begin
                    if (dataCtrl_io_stride) begin
                      if (_T_626) begin
                        state <= 3'h5;
                      end else begin
                        if (_T_618) begin
                          state <= 3'h2;
                        end else begin
                          state <= 3'h3;
                        end
                      end
                    end else begin
                      if (dataCtrl_io_split) begin
                        state <= 3'h3;
                      end
                    end
                  end
                end
              end else begin
                if (_T_633) begin
                  if (xPadCtrl1_io_done) begin
                    if (dataCtrlDone) begin
                      if (_T_628) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end else begin
                      if (_T_618) begin
                        state <= 3'h2;
                      end else begin
                        state <= 3'h3;
                      end
                    end
                  end
                end else begin
                  if (_T_638) begin
                    if (_T_639) begin
                      state <= 3'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    waddr_cur <= _GEN_37[10:0];
    waddr_nxt <= _GEN_38[10:0];
    rvalid <= io_tensor_rd_idx_valid;
    if (_GEN_51) begin
      tensorFile_0_0_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_51) begin
      tensorFile_0_1_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
  end
endmodule
module TensorDataCtrl_1( // @[:@2432.2]
  input          clock, // @[:@2433.4]
  input          io_start, // @[:@2435.4]
  output         io_done, // @[:@2435.4]
  input  [127:0] io_inst, // @[:@2435.4]
  input  [31:0]  io_baddr, // @[:@2435.4]
  input          io_xinit, // @[:@2435.4]
  input          io_xupdate, // @[:@2435.4]
  input          io_yupdate, // @[:@2435.4]
  output         io_stride, // @[:@2435.4]
  output         io_split, // @[:@2435.4]
  output [31:0]  io_addr, // @[:@2435.4]
  output [7:0]   io_len // @[:@2435.4]
);
  wire [31:0] dec_dram_offset; // @[TensorUtil.scala 251:29:@2454.4]
  wire [15:0] dec_ysize; // @[TensorUtil.scala 251:29:@2458.4]
  wire [15:0] dec_xsize; // @[TensorUtil.scala 251:29:@2460.4]
  wire [15:0] dec_xstride; // @[TensorUtil.scala 251:29:@2462.4]
  reg [31:0] caddr; // @[TensorUtil.scala 253:18:@2472.4]
  reg [31:0] _RAND_0;
  reg [31:0] baddr; // @[TensorUtil.scala 254:18:@2473.4]
  reg [31:0] _RAND_1;
  reg [7:0] len; // @[TensorUtil.scala 255:16:@2474.4]
  reg [31:0] _RAND_2;
  reg [7:0] xcnt; // @[TensorUtil.scala 267:17:@2539.4]
  reg [31:0] _RAND_3;
  reg [15:0] xrem; // @[TensorUtil.scala 268:17:@2540.4]
  reg [31:0] _RAND_4;
  wire [20:0] _GEN_27; // @[TensorUtil.scala 269:26:@2541.4]
  wire [20:0] _T_154; // @[TensorUtil.scala 269:26:@2541.4]
  wire [21:0] _T_156; // @[TensorUtil.scala 269:51:@2542.4]
  wire [21:0] _T_157; // @[TensorUtil.scala 269:51:@2543.4]
  wire [20:0] xsize; // @[TensorUtil.scala 269:51:@2544.4]
  reg [15:0] ycnt; // @[TensorUtil.scala 271:17:@2545.4]
  reg [31:0] _RAND_5;
  reg [31:0] xfer_bytes; // @[TensorUtil.scala 273:23:@2546.4]
  reg [31:0] _RAND_6;
  wire [23:0] _GEN_28; // @[TensorUtil.scala 275:35:@2547.4]
  wire [23:0] xstride_bytes; // @[TensorUtil.scala 275:35:@2547.4]
  wire [39:0] _GEN_29; // @[TensorUtil.scala 277:66:@2548.4]
  wire [39:0] _T_160; // @[TensorUtil.scala 277:66:@2548.4]
  wire [39:0] _T_161; // @[TensorUtil.scala 277:47:@2549.4]
  wire [39:0] _GEN_30; // @[TensorUtil.scala 277:33:@2550.4]
  wire [39:0] xfer_init_addr; // @[TensorUtil.scala 277:33:@2550.4]
  wire [32:0] _T_162; // @[TensorUtil.scala 278:31:@2551.4]
  wire [31:0] xfer_split_addr; // @[TensorUtil.scala 278:31:@2552.4]
  wire [31:0] _GEN_31; // @[TensorUtil.scala 279:32:@2553.4]
  wire [32:0] _T_163; // @[TensorUtil.scala 279:32:@2553.4]
  wire [31:0] xfer_stride_addr; // @[TensorUtil.scala 279:32:@2554.4]
  wire [39:0] _GEN_12; // @[TensorUtil.scala 281:55:@2555.4]
  wire [11:0] _T_164; // @[TensorUtil.scala 281:55:@2555.4]
  wire [12:0] _T_165; // @[TensorUtil.scala 281:38:@2556.4]
  wire [12:0] _T_166; // @[TensorUtil.scala 281:38:@2557.4]
  wire [11:0] xfer_init_bytes; // @[TensorUtil.scala 281:38:@2558.4]
  wire [8:0] xfer_init_pulses; // @[TensorUtil.scala 282:43:@2559.4]
  wire [31:0] _GEN_16; // @[TensorUtil.scala 283:56:@2560.4]
  wire [11:0] _T_167; // @[TensorUtil.scala 283:56:@2560.4]
  wire [12:0] _T_168; // @[TensorUtil.scala 283:38:@2561.4]
  wire [12:0] _T_169; // @[TensorUtil.scala 283:38:@2562.4]
  wire [11:0] xfer_split_bytes; // @[TensorUtil.scala 283:38:@2563.4]
  wire [8:0] xfer_split_pulses; // @[TensorUtil.scala 284:44:@2564.4]
  wire [31:0] _GEN_18; // @[TensorUtil.scala 285:57:@2565.4]
  wire [11:0] _T_170; // @[TensorUtil.scala 285:57:@2565.4]
  wire [12:0] _T_171; // @[TensorUtil.scala 285:38:@2566.4]
  wire [12:0] _T_172; // @[TensorUtil.scala 285:38:@2567.4]
  wire [11:0] xfer_stride_bytes; // @[TensorUtil.scala 285:38:@2568.4]
  wire [8:0] xfer_stride_pulses; // @[TensorUtil.scala 286:45:@2569.4]
  wire  _T_173; // @[TensorUtil.scala 288:21:@2570.4]
  wire  _T_175; // @[TensorUtil.scala 289:10:@2571.4]
  wire  _T_176; // @[TensorUtil.scala 288:29:@2572.4]
  wire [16:0] _T_178; // @[TensorUtil.scala 290:24:@2573.4]
  wire [16:0] _T_179; // @[TensorUtil.scala 290:24:@2574.4]
  wire [15:0] _T_180; // @[TensorUtil.scala 290:24:@2575.4]
  wire  _T_181; // @[TensorUtil.scala 290:10:@2576.4]
  wire  stride; // @[TensorUtil.scala 289:18:@2577.4]
  wire  _T_184; // @[TensorUtil.scala 292:35:@2579.4]
  wire  split; // @[TensorUtil.scala 292:28:@2580.4]
  wire [20:0] _GEN_32; // @[TensorUtil.scala 296:16:@2583.6]
  wire  _T_185; // @[TensorUtil.scala 296:16:@2583.6]
  wire [9:0] _T_188; // @[TensorUtil.scala 300:31:@2589.8]
  wire [9:0] _T_189; // @[TensorUtil.scala 300:31:@2590.8]
  wire [8:0] _T_190; // @[TensorUtil.scala 300:31:@2591.8]
  wire [21:0] _T_191; // @[TensorUtil.scala 301:21:@2593.8]
  wire [21:0] _T_192; // @[TensorUtil.scala 301:21:@2594.8]
  wire [20:0] _T_193; // @[TensorUtil.scala 301:21:@2595.8]
  wire [20:0] _GEN_0; // @[TensorUtil.scala 296:36:@2584.6]
  wire [20:0] _GEN_1; // @[TensorUtil.scala 296:36:@2584.6]
  wire  _T_194; // @[TensorUtil.scala 303:25:@2600.6]
  wire [20:0] _GEN_34; // @[TensorUtil.scala 305:16:@2603.8]
  wire  _T_195; // @[TensorUtil.scala 305:16:@2603.8]
  wire [9:0] _T_198; // @[TensorUtil.scala 309:33:@2609.10]
  wire [9:0] _T_199; // @[TensorUtil.scala 309:33:@2610.10]
  wire [8:0] _T_200; // @[TensorUtil.scala 309:33:@2611.10]
  wire [21:0] _T_201; // @[TensorUtil.scala 310:21:@2613.10]
  wire [21:0] _T_202; // @[TensorUtil.scala 310:21:@2614.10]
  wire [20:0] _T_203; // @[TensorUtil.scala 310:21:@2615.10]
  wire [20:0] _GEN_2; // @[TensorUtil.scala 305:38:@2604.8]
  wire [20:0] _GEN_3; // @[TensorUtil.scala 305:38:@2604.8]
  wire  _T_204; // @[TensorUtil.scala 312:25:@2620.8]
  wire [15:0] _GEN_36; // @[TensorUtil.scala 314:15:@2623.10]
  wire  _T_205; // @[TensorUtil.scala 314:15:@2623.10]
  wire [9:0] _T_208; // @[TensorUtil.scala 318:32:@2629.12]
  wire [9:0] _T_209; // @[TensorUtil.scala 318:32:@2630.12]
  wire [8:0] _T_210; // @[TensorUtil.scala 318:32:@2631.12]
  wire [16:0] _T_211; // @[TensorUtil.scala 319:20:@2633.12]
  wire [16:0] _T_212; // @[TensorUtil.scala 319:20:@2634.12]
  wire [15:0] _T_213; // @[TensorUtil.scala 319:20:@2635.12]
  wire [15:0] _GEN_4; // @[TensorUtil.scala 314:36:@2624.10]
  wire [15:0] _GEN_5; // @[TensorUtil.scala 314:36:@2624.10]
  wire [31:0] _GEN_6; // @[TensorUtil.scala 312:35:@2621.8]
  wire [15:0] _GEN_7; // @[TensorUtil.scala 312:35:@2621.8]
  wire [15:0] _GEN_8; // @[TensorUtil.scala 312:35:@2621.8]
  wire [31:0] _GEN_9; // @[TensorUtil.scala 303:36:@2601.6]
  wire [20:0] _GEN_10; // @[TensorUtil.scala 303:36:@2601.6]
  wire [20:0] _GEN_11; // @[TensorUtil.scala 303:36:@2601.6]
  wire [20:0] _GEN_13; // @[TensorUtil.scala 294:18:@2581.4]
  wire [20:0] _GEN_14; // @[TensorUtil.scala 294:18:@2581.4]
  wire [8:0] _T_216; // @[TensorUtil.scala 326:18:@2644.8]
  wire [7:0] _T_217; // @[TensorUtil.scala 326:18:@2645.8]
  wire [7:0] _GEN_15; // @[TensorUtil.scala 325:26:@2643.6]
  wire  _T_219; // @[TensorUtil.scala 331:25:@2652.6]
  wire [16:0] _T_221; // @[TensorUtil.scala 332:18:@2654.8]
  wire [15:0] _T_222; // @[TensorUtil.scala 332:18:@2655.8]
  wire [15:0] _GEN_17; // @[TensorUtil.scala 331:36:@2653.6]
  wire [31:0] _GEN_19; // @[TensorUtil.scala 341:24:@2668.10]
  wire [31:0] _GEN_20; // @[TensorUtil.scala 341:24:@2668.10]
  wire [31:0] _GEN_21; // @[TensorUtil.scala 339:17:@2664.8]
  wire [31:0] _GEN_22; // @[TensorUtil.scala 339:17:@2664.8]
  wire [31:0] _GEN_23; // @[TensorUtil.scala 338:26:@2663.6]
  wire [31:0] _GEN_24; // @[TensorUtil.scala 338:26:@2663.6]
  wire [39:0] _GEN_25; // @[TensorUtil.scala 335:18:@2658.4]
  wire [39:0] _GEN_26; // @[TensorUtil.scala 335:18:@2658.4]
  wire  _T_232; // @[TensorUtil.scala 354:10:@2685.4]
  assign dec_dram_offset = io_inst[56:25]; // @[TensorUtil.scala 251:29:@2454.4]
  assign dec_ysize = io_inst[79:64]; // @[TensorUtil.scala 251:29:@2458.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 251:29:@2460.4]
  assign dec_xstride = io_inst[111:96]; // @[TensorUtil.scala 251:29:@2462.4]
  assign _GEN_27 = {{5'd0}, dec_xsize}; // @[TensorUtil.scala 269:26:@2541.4]
  assign _T_154 = _GEN_27 << 5; // @[TensorUtil.scala 269:26:@2541.4]
  assign _T_156 = _T_154 - 21'h1; // @[TensorUtil.scala 269:51:@2542.4]
  assign _T_157 = $unsigned(_T_156); // @[TensorUtil.scala 269:51:@2543.4]
  assign xsize = _T_157[20:0]; // @[TensorUtil.scala 269:51:@2544.4]
  assign _GEN_28 = {{8'd0}, dec_xstride}; // @[TensorUtil.scala 275:35:@2547.4]
  assign xstride_bytes = _GEN_28 << 8; // @[TensorUtil.scala 275:35:@2547.4]
  assign _GEN_29 = {{8'd0}, dec_dram_offset}; // @[TensorUtil.scala 277:66:@2548.4]
  assign _T_160 = _GEN_29 << 8; // @[TensorUtil.scala 277:66:@2548.4]
  assign _T_161 = 40'hffffffff & _T_160; // @[TensorUtil.scala 277:47:@2549.4]
  assign _GEN_30 = {{8'd0}, io_baddr}; // @[TensorUtil.scala 277:33:@2550.4]
  assign xfer_init_addr = _GEN_30 | _T_161; // @[TensorUtil.scala 277:33:@2550.4]
  assign _T_162 = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@2551.4]
  assign xfer_split_addr = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@2552.4]
  assign _GEN_31 = {{8'd0}, xstride_bytes}; // @[TensorUtil.scala 279:32:@2553.4]
  assign _T_163 = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@2553.4]
  assign xfer_stride_addr = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@2554.4]
  assign _GEN_12 = xfer_init_addr % 40'h800; // @[TensorUtil.scala 281:55:@2555.4]
  assign _T_164 = _GEN_12[11:0]; // @[TensorUtil.scala 281:55:@2555.4]
  assign _T_165 = 12'h800 - _T_164; // @[TensorUtil.scala 281:38:@2556.4]
  assign _T_166 = $unsigned(_T_165); // @[TensorUtil.scala 281:38:@2557.4]
  assign xfer_init_bytes = _T_166[11:0]; // @[TensorUtil.scala 281:38:@2558.4]
  assign xfer_init_pulses = xfer_init_bytes[11:3]; // @[TensorUtil.scala 282:43:@2559.4]
  assign _GEN_16 = xfer_split_addr % 32'h800; // @[TensorUtil.scala 283:56:@2560.4]
  assign _T_167 = _GEN_16[11:0]; // @[TensorUtil.scala 283:56:@2560.4]
  assign _T_168 = 12'h800 - _T_167; // @[TensorUtil.scala 283:38:@2561.4]
  assign _T_169 = $unsigned(_T_168); // @[TensorUtil.scala 283:38:@2562.4]
  assign xfer_split_bytes = _T_169[11:0]; // @[TensorUtil.scala 283:38:@2563.4]
  assign xfer_split_pulses = xfer_split_bytes[11:3]; // @[TensorUtil.scala 284:44:@2564.4]
  assign _GEN_18 = xfer_stride_addr % 32'h800; // @[TensorUtil.scala 285:57:@2565.4]
  assign _T_170 = _GEN_18[11:0]; // @[TensorUtil.scala 285:57:@2565.4]
  assign _T_171 = 12'h800 - _T_170; // @[TensorUtil.scala 285:38:@2566.4]
  assign _T_172 = $unsigned(_T_171); // @[TensorUtil.scala 285:38:@2567.4]
  assign xfer_stride_bytes = _T_172[11:0]; // @[TensorUtil.scala 285:38:@2568.4]
  assign xfer_stride_pulses = xfer_stride_bytes[11:3]; // @[TensorUtil.scala 286:45:@2569.4]
  assign _T_173 = xcnt == len; // @[TensorUtil.scala 288:21:@2570.4]
  assign _T_175 = xrem == 16'h0; // @[TensorUtil.scala 289:10:@2571.4]
  assign _T_176 = _T_173 & _T_175; // @[TensorUtil.scala 288:29:@2572.4]
  assign _T_178 = dec_ysize - 16'h1; // @[TensorUtil.scala 290:24:@2573.4]
  assign _T_179 = $unsigned(_T_178); // @[TensorUtil.scala 290:24:@2574.4]
  assign _T_180 = _T_179[15:0]; // @[TensorUtil.scala 290:24:@2575.4]
  assign _T_181 = ycnt != _T_180; // @[TensorUtil.scala 290:10:@2576.4]
  assign stride = _T_176 & _T_181; // @[TensorUtil.scala 289:18:@2577.4]
  assign _T_184 = xrem != 16'h0; // @[TensorUtil.scala 292:35:@2579.4]
  assign split = _T_173 & _T_184; // @[TensorUtil.scala 292:28:@2580.4]
  assign _GEN_32 = {{12'd0}, xfer_init_pulses}; // @[TensorUtil.scala 296:16:@2583.6]
  assign _T_185 = xsize < _GEN_32; // @[TensorUtil.scala 296:16:@2583.6]
  assign _T_188 = xfer_init_pulses - 9'h1; // @[TensorUtil.scala 300:31:@2589.8]
  assign _T_189 = $unsigned(_T_188); // @[TensorUtil.scala 300:31:@2590.8]
  assign _T_190 = _T_189[8:0]; // @[TensorUtil.scala 300:31:@2591.8]
  assign _T_191 = xsize - _GEN_32; // @[TensorUtil.scala 301:21:@2593.8]
  assign _T_192 = $unsigned(_T_191); // @[TensorUtil.scala 301:21:@2594.8]
  assign _T_193 = _T_192[20:0]; // @[TensorUtil.scala 301:21:@2595.8]
  assign _GEN_0 = _T_185 ? xsize : {{12'd0}, _T_190}; // @[TensorUtil.scala 296:36:@2584.6]
  assign _GEN_1 = _T_185 ? 21'h0 : _T_193; // @[TensorUtil.scala 296:36:@2584.6]
  assign _T_194 = io_xupdate & stride; // @[TensorUtil.scala 303:25:@2600.6]
  assign _GEN_34 = {{12'd0}, xfer_stride_pulses}; // @[TensorUtil.scala 305:16:@2603.8]
  assign _T_195 = xsize < _GEN_34; // @[TensorUtil.scala 305:16:@2603.8]
  assign _T_198 = xfer_stride_pulses - 9'h1; // @[TensorUtil.scala 309:33:@2609.10]
  assign _T_199 = $unsigned(_T_198); // @[TensorUtil.scala 309:33:@2610.10]
  assign _T_200 = _T_199[8:0]; // @[TensorUtil.scala 309:33:@2611.10]
  assign _T_201 = xsize - _GEN_34; // @[TensorUtil.scala 310:21:@2613.10]
  assign _T_202 = $unsigned(_T_201); // @[TensorUtil.scala 310:21:@2614.10]
  assign _T_203 = _T_202[20:0]; // @[TensorUtil.scala 310:21:@2615.10]
  assign _GEN_2 = _T_195 ? xsize : {{12'd0}, _T_200}; // @[TensorUtil.scala 305:38:@2604.8]
  assign _GEN_3 = _T_195 ? 21'h0 : _T_203; // @[TensorUtil.scala 305:38:@2604.8]
  assign _T_204 = io_xupdate & split; // @[TensorUtil.scala 312:25:@2620.8]
  assign _GEN_36 = {{7'd0}, xfer_split_pulses}; // @[TensorUtil.scala 314:15:@2623.10]
  assign _T_205 = xrem < _GEN_36; // @[TensorUtil.scala 314:15:@2623.10]
  assign _T_208 = xfer_split_pulses - 9'h1; // @[TensorUtil.scala 318:32:@2629.12]
  assign _T_209 = $unsigned(_T_208); // @[TensorUtil.scala 318:32:@2630.12]
  assign _T_210 = _T_209[8:0]; // @[TensorUtil.scala 318:32:@2631.12]
  assign _T_211 = xrem - _GEN_36; // @[TensorUtil.scala 319:20:@2633.12]
  assign _T_212 = $unsigned(_T_211); // @[TensorUtil.scala 319:20:@2634.12]
  assign _T_213 = _T_212[15:0]; // @[TensorUtil.scala 319:20:@2635.12]
  assign _GEN_4 = _T_205 ? xrem : {{7'd0}, _T_210}; // @[TensorUtil.scala 314:36:@2624.10]
  assign _GEN_5 = _T_205 ? 16'h0 : _T_213; // @[TensorUtil.scala 314:36:@2624.10]
  assign _GEN_6 = _T_204 ? {{20'd0}, xfer_split_bytes} : xfer_bytes; // @[TensorUtil.scala 312:35:@2621.8]
  assign _GEN_7 = _T_204 ? _GEN_4 : {{8'd0}, len}; // @[TensorUtil.scala 312:35:@2621.8]
  assign _GEN_8 = _T_204 ? _GEN_5 : xrem; // @[TensorUtil.scala 312:35:@2621.8]
  assign _GEN_9 = _T_194 ? {{20'd0}, xfer_stride_bytes} : _GEN_6; // @[TensorUtil.scala 303:36:@2601.6]
  assign _GEN_10 = _T_194 ? _GEN_2 : {{5'd0}, _GEN_7}; // @[TensorUtil.scala 303:36:@2601.6]
  assign _GEN_11 = _T_194 ? _GEN_3 : {{5'd0}, _GEN_8}; // @[TensorUtil.scala 303:36:@2601.6]
  assign _GEN_13 = io_start ? _GEN_0 : _GEN_10; // @[TensorUtil.scala 294:18:@2581.4]
  assign _GEN_14 = io_start ? _GEN_1 : _GEN_11; // @[TensorUtil.scala 294:18:@2581.4]
  assign _T_216 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@2644.8]
  assign _T_217 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@2645.8]
  assign _GEN_15 = io_xupdate ? _T_217 : xcnt; // @[TensorUtil.scala 325:26:@2643.6]
  assign _T_219 = io_yupdate & stride; // @[TensorUtil.scala 331:25:@2652.6]
  assign _T_221 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@2654.8]
  assign _T_222 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@2655.8]
  assign _GEN_17 = _T_219 ? _T_222 : ycnt; // @[TensorUtil.scala 331:36:@2653.6]
  assign _GEN_19 = stride ? xfer_stride_addr : caddr; // @[TensorUtil.scala 341:24:@2668.10]
  assign _GEN_20 = stride ? xfer_stride_addr : baddr; // @[TensorUtil.scala 341:24:@2668.10]
  assign _GEN_21 = split ? xfer_split_addr : _GEN_19; // @[TensorUtil.scala 339:17:@2664.8]
  assign _GEN_22 = split ? baddr : _GEN_20; // @[TensorUtil.scala 339:17:@2664.8]
  assign _GEN_23 = io_yupdate ? _GEN_21 : caddr; // @[TensorUtil.scala 338:26:@2663.6]
  assign _GEN_24 = io_yupdate ? _GEN_22 : baddr; // @[TensorUtil.scala 338:26:@2663.6]
  assign _GEN_25 = io_start ? xfer_init_addr : {{8'd0}, _GEN_23}; // @[TensorUtil.scala 335:18:@2658.4]
  assign _GEN_26 = io_start ? xfer_init_addr : {{8'd0}, _GEN_24}; // @[TensorUtil.scala 335:18:@2658.4]
  assign _T_232 = ycnt == _T_180; // @[TensorUtil.scala 354:10:@2685.4]
  assign io_done = _T_176 & _T_232; // @[TensorUtil.scala 352:11:@2687.4]
  assign io_stride = _T_176 & _T_181; // @[TensorUtil.scala 347:13:@2673.4]
  assign io_split = _T_173 & _T_184; // @[TensorUtil.scala 348:12:@2674.4]
  assign io_addr = caddr; // @[TensorUtil.scala 350:11:@2677.4]
  assign io_len = len; // @[TensorUtil.scala 351:10:@2678.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  caddr = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  baddr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  len = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  xcnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xrem = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ycnt = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  xfer_bytes = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    caddr <= _GEN_25[31:0];
    baddr <= _GEN_26[31:0];
    len <= _GEN_13[7:0];
    if (io_xinit) begin
      xcnt <= 8'h0;
    end else begin
      if (io_xupdate) begin
        xcnt <= _T_217;
      end
    end
    xrem <= _GEN_14[15:0];
    if (io_start) begin
      ycnt <= 16'h0;
    end else begin
      if (_T_219) begin
        ycnt <= _T_222;
      end
    end
    if (io_start) begin
      xfer_bytes <= {{20'd0}, xfer_init_bytes};
    end else begin
      if (_T_194) begin
        xfer_bytes <= {{20'd0}, xfer_stride_bytes};
      end else begin
        if (_T_204) begin
          xfer_bytes <= {{20'd0}, xfer_split_bytes};
        end
      end
    end
  end
endmodule
module TensorPadCtrl_4( // @[:@2689.2]
  input          clock, // @[:@2690.4]
  input          reset, // @[:@2691.4]
  input          io_start, // @[:@2692.4]
  output         io_done, // @[:@2692.4]
  input  [127:0] io_inst // @[:@2692.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@2717.4]
  wire [3:0] dec_ypad_0; // @[TensorUtil.scala 173:29:@2721.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@2725.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@2727.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@2729.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@2730.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@2731.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@2732.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@2733.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@2733.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@2734.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@2735.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@2735.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@2736.4]
  wire [20:0] _GEN_12; // @[TensorUtil.scala 182:46:@2737.4]
  wire [20:0] _T_39; // @[TensorUtil.scala 182:46:@2737.4]
  wire [21:0] _T_41; // @[TensorUtil.scala 182:71:@2738.4]
  wire [21:0] _T_42; // @[TensorUtil.scala 182:71:@2739.4]
  wire [20:0] xval; // @[TensorUtil.scala 182:71:@2740.4]
  wire  _T_44; // @[TensorUtil.scala 190:22:@2741.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 190:42:@2742.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 190:42:@2743.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 190:42:@2744.4]
  wire [3:0] yval; // @[TensorUtil.scala 190:10:@2745.4]
  reg  state; // @[TensorUtil.scala 197:22:@2746.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@2747.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@2749.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@2756.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@2757.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@2758.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@2759.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@2755.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@2748.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@2763.4]
  wire [20:0] _GEN_4; // @[TensorUtil.scala 212:25:@2764.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@2770.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@2777.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@2778.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@2776.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@2782.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@2783.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@2790.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@2792.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@2793.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@2791.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@2798.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@2717.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorUtil.scala 173:29:@2721.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@2725.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@2727.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@2733.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@2733.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@2734.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@2735.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@2735.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@2736.4]
  assign _GEN_12 = {{5'd0}, _T_38}; // @[TensorUtil.scala 182:46:@2737.4]
  assign _T_39 = _GEN_12 << 5; // @[TensorUtil.scala 182:46:@2737.4]
  assign _T_41 = _T_39 - 21'h1; // @[TensorUtil.scala 182:71:@2738.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@2739.4]
  assign xval = _T_42[20:0]; // @[TensorUtil.scala 182:71:@2740.4]
  assign _T_44 = dec_ypad_0 != 4'h0; // @[TensorUtil.scala 190:22:@2741.4]
  assign _T_46 = dec_ypad_0 - 4'h1; // @[TensorUtil.scala 190:42:@2742.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 190:42:@2743.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 190:42:@2744.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 190:10:@2745.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@2747.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@2749.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@2756.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@2757.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@2758.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@2759.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@2755.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@2748.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@2763.4]
  assign _GEN_4 = _T_56 ? xval : {{5'd0}, xmax}; // @[TensorUtil.scala 212:25:@2764.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@2770.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2777.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2778.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@2776.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@2782.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@2783.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@2790.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@2792.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@2793.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@2791.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@2798.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@2801.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_5( // @[:@2803.2]
  input          clock, // @[:@2804.4]
  input          reset, // @[:@2805.4]
  input          io_start, // @[:@2806.4]
  output         io_done, // @[:@2806.4]
  input  [127:0] io_inst // @[:@2806.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@2831.4]
  wire [3:0] dec_ypad_1; // @[TensorUtil.scala 173:29:@2837.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@2839.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@2841.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@2843.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@2844.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@2845.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@2846.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@2847.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@2847.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@2848.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@2849.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@2849.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@2850.4]
  wire [20:0] _GEN_12; // @[TensorUtil.scala 182:46:@2851.4]
  wire [20:0] _T_39; // @[TensorUtil.scala 182:46:@2851.4]
  wire [21:0] _T_41; // @[TensorUtil.scala 182:71:@2852.4]
  wire [21:0] _T_42; // @[TensorUtil.scala 182:71:@2853.4]
  wire [20:0] xval; // @[TensorUtil.scala 182:71:@2854.4]
  wire  _T_44; // @[TensorUtil.scala 192:22:@2855.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 192:42:@2856.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 192:42:@2857.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 192:42:@2858.4]
  wire [3:0] yval; // @[TensorUtil.scala 192:10:@2859.4]
  reg  state; // @[TensorUtil.scala 197:22:@2860.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@2861.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@2863.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@2870.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@2871.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@2872.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@2873.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@2869.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@2862.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@2877.4]
  wire [20:0] _GEN_4; // @[TensorUtil.scala 212:25:@2878.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@2884.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@2891.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@2892.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@2890.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@2896.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@2897.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@2904.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@2906.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@2907.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@2905.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@2912.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@2831.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorUtil.scala 173:29:@2837.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@2839.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@2841.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@2847.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@2847.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@2848.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@2849.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@2849.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@2850.4]
  assign _GEN_12 = {{5'd0}, _T_38}; // @[TensorUtil.scala 182:46:@2851.4]
  assign _T_39 = _GEN_12 << 5; // @[TensorUtil.scala 182:46:@2851.4]
  assign _T_41 = _T_39 - 21'h1; // @[TensorUtil.scala 182:71:@2852.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@2853.4]
  assign xval = _T_42[20:0]; // @[TensorUtil.scala 182:71:@2854.4]
  assign _T_44 = dec_ypad_1 != 4'h0; // @[TensorUtil.scala 192:22:@2855.4]
  assign _T_46 = dec_ypad_1 - 4'h1; // @[TensorUtil.scala 192:42:@2856.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 192:42:@2857.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 192:42:@2858.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 192:10:@2859.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@2861.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@2863.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@2870.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@2871.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@2872.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@2873.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@2869.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@2862.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@2877.4]
  assign _GEN_4 = _T_56 ? xval : {{5'd0}, xmax}; // @[TensorUtil.scala 212:25:@2878.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@2884.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2891.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2892.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@2890.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@2896.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@2897.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@2904.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@2906.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@2907.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@2905.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@2912.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@2915.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_6( // @[:@2917.2]
  input          clock, // @[:@2918.4]
  input          reset, // @[:@2919.4]
  input          io_start, // @[:@2920.4]
  output         io_done, // @[:@2920.4]
  input  [127:0] io_inst // @[:@2920.4]
);
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@2953.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@2957.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@2959.4]
  reg [31:0] _RAND_1;
  wire [8:0] _GEN_10; // @[TensorUtil.scala 184:19:@2961.4]
  wire [8:0] _T_35; // @[TensorUtil.scala 184:19:@2961.4]
  wire [9:0] _T_37; // @[TensorUtil.scala 184:44:@2962.4]
  wire [9:0] _T_38; // @[TensorUtil.scala 184:44:@2963.4]
  wire [8:0] xval; // @[TensorUtil.scala 184:44:@2964.4]
  reg  state; // @[TensorUtil.scala 197:22:@2965.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@2966.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@2968.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@2976.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@2978.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@2974.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@2967.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@2982.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@2989.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@2996.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@2997.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@2995.6]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@2953.4]
  assign _GEN_10 = {{5'd0}, dec_xpad_0}; // @[TensorUtil.scala 184:19:@2961.4]
  assign _T_35 = _GEN_10 << 5; // @[TensorUtil.scala 184:19:@2961.4]
  assign _T_37 = _T_35 - 9'h1; // @[TensorUtil.scala 184:44:@2962.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 184:44:@2963.4]
  assign xval = _T_38[8:0]; // @[TensorUtil.scala 184:44:@2964.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@2966.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@2968.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@2976.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@2978.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@2974.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@2967.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@2982.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@2989.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2996.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@2997.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@2995.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@3020.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{7'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_7( // @[:@3022.2]
  input          clock, // @[:@3023.4]
  input          reset, // @[:@3024.4]
  input          io_start, // @[:@3025.4]
  output         io_done, // @[:@3025.4]
  input  [127:0] io_inst // @[:@3025.4]
);
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@3060.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@3062.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@3064.4]
  reg [31:0] _RAND_1;
  wire [8:0] _GEN_10; // @[TensorUtil.scala 186:19:@3066.4]
  wire [8:0] _T_35; // @[TensorUtil.scala 186:19:@3066.4]
  wire [9:0] _T_37; // @[TensorUtil.scala 186:44:@3067.4]
  wire [9:0] _T_38; // @[TensorUtil.scala 186:44:@3068.4]
  wire [8:0] xval; // @[TensorUtil.scala 186:44:@3069.4]
  reg  state; // @[TensorUtil.scala 197:22:@3070.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@3071.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@3073.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@3081.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@3083.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@3079.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@3072.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@3087.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@3094.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@3101.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@3102.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@3100.6]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@3060.4]
  assign _GEN_10 = {{5'd0}, dec_xpad_1}; // @[TensorUtil.scala 186:19:@3066.4]
  assign _T_35 = _GEN_10 << 5; // @[TensorUtil.scala 186:19:@3066.4]
  assign _T_37 = _T_35 - 9'h1; // @[TensorUtil.scala 186:44:@3067.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 186:44:@3068.4]
  assign xval = _T_38[8:0]; // @[TensorUtil.scala 186:44:@3069.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@3071.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@3073.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@3081.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@3083.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@3079.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@3072.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@3087.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@3094.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@3101.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@3102.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@3100.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@3125.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{7'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorLoad_1( // @[:@3127.2]
  input          clock, // @[:@3128.4]
  input          reset, // @[:@3129.4]
  input          io_start, // @[:@3130.4]
  output         io_done, // @[:@3130.4]
  input  [127:0] io_inst, // @[:@3130.4]
  input  [31:0]  io_baddr, // @[:@3130.4]
  input          io_vme_rd_cmd_ready, // @[:@3130.4]
  output         io_vme_rd_cmd_valid, // @[:@3130.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@3130.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@3130.4]
  output         io_vme_rd_data_ready, // @[:@3130.4]
  input          io_vme_rd_data_valid, // @[:@3130.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@3130.4]
  input          io_tensor_rd_idx_valid, // @[:@3130.4]
  input  [9:0]   io_tensor_rd_idx_bits, // @[:@3130.4]
  output         io_tensor_rd_data_valid, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_0_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_1_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_2_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_3_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_4_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_5_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_6_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_7_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_8_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_9_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_10_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_11_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_12_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_13_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_14_15, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_0, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_1, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_2, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_3, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_4, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_5, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_6, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_7, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_8, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_9, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_10, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_11, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_12, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_13, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_14, // @[:@3130.4]
  output [7:0]   io_tensor_rd_data_bits_15_15 // @[:@3130.4]
);
  wire  dataCtrl_clock; // @[TensorLoad.scala 52:24:@3167.4]
  wire  dataCtrl_io_start; // @[TensorLoad.scala 52:24:@3167.4]
  wire  dataCtrl_io_done; // @[TensorLoad.scala 52:24:@3167.4]
  wire [127:0] dataCtrl_io_inst; // @[TensorLoad.scala 52:24:@3167.4]
  wire [31:0] dataCtrl_io_baddr; // @[TensorLoad.scala 52:24:@3167.4]
  wire  dataCtrl_io_xinit; // @[TensorLoad.scala 52:24:@3167.4]
  wire  dataCtrl_io_xupdate; // @[TensorLoad.scala 52:24:@3167.4]
  wire  dataCtrl_io_yupdate; // @[TensorLoad.scala 52:24:@3167.4]
  wire  dataCtrl_io_stride; // @[TensorLoad.scala 52:24:@3167.4]
  wire  dataCtrl_io_split; // @[TensorLoad.scala 52:24:@3167.4]
  wire [31:0] dataCtrl_io_addr; // @[TensorLoad.scala 52:24:@3167.4]
  wire [7:0] dataCtrl_io_len; // @[TensorLoad.scala 52:24:@3167.4]
  wire  yPadCtrl0_clock; // @[TensorLoad.scala 55:25:@3171.4]
  wire  yPadCtrl0_reset; // @[TensorLoad.scala 55:25:@3171.4]
  wire  yPadCtrl0_io_start; // @[TensorLoad.scala 55:25:@3171.4]
  wire  yPadCtrl0_io_done; // @[TensorLoad.scala 55:25:@3171.4]
  wire [127:0] yPadCtrl0_io_inst; // @[TensorLoad.scala 55:25:@3171.4]
  wire  yPadCtrl1_clock; // @[TensorLoad.scala 56:25:@3174.4]
  wire  yPadCtrl1_reset; // @[TensorLoad.scala 56:25:@3174.4]
  wire  yPadCtrl1_io_start; // @[TensorLoad.scala 56:25:@3174.4]
  wire  yPadCtrl1_io_done; // @[TensorLoad.scala 56:25:@3174.4]
  wire [127:0] yPadCtrl1_io_inst; // @[TensorLoad.scala 56:25:@3174.4]
  wire  xPadCtrl0_clock; // @[TensorLoad.scala 57:25:@3177.4]
  wire  xPadCtrl0_reset; // @[TensorLoad.scala 57:25:@3177.4]
  wire  xPadCtrl0_io_start; // @[TensorLoad.scala 57:25:@3177.4]
  wire  xPadCtrl0_io_done; // @[TensorLoad.scala 57:25:@3177.4]
  wire [127:0] xPadCtrl0_io_inst; // @[TensorLoad.scala 57:25:@3177.4]
  wire  xPadCtrl1_clock; // @[TensorLoad.scala 58:25:@3180.4]
  wire  xPadCtrl1_reset; // @[TensorLoad.scala 58:25:@3180.4]
  wire  xPadCtrl1_io_start; // @[TensorLoad.scala 58:25:@3180.4]
  wire  xPadCtrl1_io_done; // @[TensorLoad.scala 58:25:@3180.4]
  wire [127:0] xPadCtrl1_io_inst; // @[TensorLoad.scala 58:25:@3180.4]
  reg [63:0] tensorFile_0_0 [0:1023]; // @[TensorLoad.scala 222:16:@3450.4]
  reg [63:0] _RAND_0;
  wire [63:0] tensorFile_0_0_rdata_0_data; // @[TensorLoad.scala 222:16:@3450.4]
  wire [9:0] tensorFile_0_0_rdata_0_addr; // @[TensorLoad.scala 222:16:@3450.4]
  wire [63:0] tensorFile_0_0__T_4976_data; // @[TensorLoad.scala 222:16:@3450.4]
  wire [9:0] tensorFile_0_0__T_4976_addr; // @[TensorLoad.scala 222:16:@3450.4]
  wire  tensorFile_0_0__T_4976_mask; // @[TensorLoad.scala 222:16:@3450.4]
  wire  tensorFile_0_0__T_4976_en; // @[TensorLoad.scala 222:16:@3450.4]
  reg [63:0] tensorFile_0_1 [0:1023]; // @[TensorLoad.scala 222:16:@3450.4]
  reg [63:0] _RAND_1;
  wire [63:0] tensorFile_0_1_rdata_0_data; // @[TensorLoad.scala 222:16:@3450.4]
  wire [9:0] tensorFile_0_1_rdata_0_addr; // @[TensorLoad.scala 222:16:@3450.4]
  wire [63:0] tensorFile_0_1__T_4976_data; // @[TensorLoad.scala 222:16:@3450.4]
  wire [9:0] tensorFile_0_1__T_4976_addr; // @[TensorLoad.scala 222:16:@3450.4]
  wire  tensorFile_0_1__T_4976_mask; // @[TensorLoad.scala 222:16:@3450.4]
  wire  tensorFile_0_1__T_4976_en; // @[TensorLoad.scala 222:16:@3450.4]
  reg [63:0] tensorFile_1_0 [0:1023]; // @[TensorLoad.scala 222:16:@3451.4]
  reg [63:0] _RAND_2;
  wire [63:0] tensorFile_1_0_rdata_1_data; // @[TensorLoad.scala 222:16:@3451.4]
  wire [9:0] tensorFile_1_0_rdata_1_addr; // @[TensorLoad.scala 222:16:@3451.4]
  wire [63:0] tensorFile_1_0__T_5063_data; // @[TensorLoad.scala 222:16:@3451.4]
  wire [9:0] tensorFile_1_0__T_5063_addr; // @[TensorLoad.scala 222:16:@3451.4]
  wire  tensorFile_1_0__T_5063_mask; // @[TensorLoad.scala 222:16:@3451.4]
  wire  tensorFile_1_0__T_5063_en; // @[TensorLoad.scala 222:16:@3451.4]
  reg [63:0] tensorFile_1_1 [0:1023]; // @[TensorLoad.scala 222:16:@3451.4]
  reg [63:0] _RAND_3;
  wire [63:0] tensorFile_1_1_rdata_1_data; // @[TensorLoad.scala 222:16:@3451.4]
  wire [9:0] tensorFile_1_1_rdata_1_addr; // @[TensorLoad.scala 222:16:@3451.4]
  wire [63:0] tensorFile_1_1__T_5063_data; // @[TensorLoad.scala 222:16:@3451.4]
  wire [9:0] tensorFile_1_1__T_5063_addr; // @[TensorLoad.scala 222:16:@3451.4]
  wire  tensorFile_1_1__T_5063_mask; // @[TensorLoad.scala 222:16:@3451.4]
  wire  tensorFile_1_1__T_5063_en; // @[TensorLoad.scala 222:16:@3451.4]
  reg [63:0] tensorFile_2_0 [0:1023]; // @[TensorLoad.scala 222:16:@3452.4]
  reg [63:0] _RAND_4;
  wire [63:0] tensorFile_2_0_rdata_2_data; // @[TensorLoad.scala 222:16:@3452.4]
  wire [9:0] tensorFile_2_0_rdata_2_addr; // @[TensorLoad.scala 222:16:@3452.4]
  wire [63:0] tensorFile_2_0__T_5150_data; // @[TensorLoad.scala 222:16:@3452.4]
  wire [9:0] tensorFile_2_0__T_5150_addr; // @[TensorLoad.scala 222:16:@3452.4]
  wire  tensorFile_2_0__T_5150_mask; // @[TensorLoad.scala 222:16:@3452.4]
  wire  tensorFile_2_0__T_5150_en; // @[TensorLoad.scala 222:16:@3452.4]
  reg [63:0] tensorFile_2_1 [0:1023]; // @[TensorLoad.scala 222:16:@3452.4]
  reg [63:0] _RAND_5;
  wire [63:0] tensorFile_2_1_rdata_2_data; // @[TensorLoad.scala 222:16:@3452.4]
  wire [9:0] tensorFile_2_1_rdata_2_addr; // @[TensorLoad.scala 222:16:@3452.4]
  wire [63:0] tensorFile_2_1__T_5150_data; // @[TensorLoad.scala 222:16:@3452.4]
  wire [9:0] tensorFile_2_1__T_5150_addr; // @[TensorLoad.scala 222:16:@3452.4]
  wire  tensorFile_2_1__T_5150_mask; // @[TensorLoad.scala 222:16:@3452.4]
  wire  tensorFile_2_1__T_5150_en; // @[TensorLoad.scala 222:16:@3452.4]
  reg [63:0] tensorFile_3_0 [0:1023]; // @[TensorLoad.scala 222:16:@3453.4]
  reg [63:0] _RAND_6;
  wire [63:0] tensorFile_3_0_rdata_3_data; // @[TensorLoad.scala 222:16:@3453.4]
  wire [9:0] tensorFile_3_0_rdata_3_addr; // @[TensorLoad.scala 222:16:@3453.4]
  wire [63:0] tensorFile_3_0__T_5237_data; // @[TensorLoad.scala 222:16:@3453.4]
  wire [9:0] tensorFile_3_0__T_5237_addr; // @[TensorLoad.scala 222:16:@3453.4]
  wire  tensorFile_3_0__T_5237_mask; // @[TensorLoad.scala 222:16:@3453.4]
  wire  tensorFile_3_0__T_5237_en; // @[TensorLoad.scala 222:16:@3453.4]
  reg [63:0] tensorFile_3_1 [0:1023]; // @[TensorLoad.scala 222:16:@3453.4]
  reg [63:0] _RAND_7;
  wire [63:0] tensorFile_3_1_rdata_3_data; // @[TensorLoad.scala 222:16:@3453.4]
  wire [9:0] tensorFile_3_1_rdata_3_addr; // @[TensorLoad.scala 222:16:@3453.4]
  wire [63:0] tensorFile_3_1__T_5237_data; // @[TensorLoad.scala 222:16:@3453.4]
  wire [9:0] tensorFile_3_1__T_5237_addr; // @[TensorLoad.scala 222:16:@3453.4]
  wire  tensorFile_3_1__T_5237_mask; // @[TensorLoad.scala 222:16:@3453.4]
  wire  tensorFile_3_1__T_5237_en; // @[TensorLoad.scala 222:16:@3453.4]
  reg [63:0] tensorFile_4_0 [0:1023]; // @[TensorLoad.scala 222:16:@3454.4]
  reg [63:0] _RAND_8;
  wire [63:0] tensorFile_4_0_rdata_4_data; // @[TensorLoad.scala 222:16:@3454.4]
  wire [9:0] tensorFile_4_0_rdata_4_addr; // @[TensorLoad.scala 222:16:@3454.4]
  wire [63:0] tensorFile_4_0__T_5324_data; // @[TensorLoad.scala 222:16:@3454.4]
  wire [9:0] tensorFile_4_0__T_5324_addr; // @[TensorLoad.scala 222:16:@3454.4]
  wire  tensorFile_4_0__T_5324_mask; // @[TensorLoad.scala 222:16:@3454.4]
  wire  tensorFile_4_0__T_5324_en; // @[TensorLoad.scala 222:16:@3454.4]
  reg [63:0] tensorFile_4_1 [0:1023]; // @[TensorLoad.scala 222:16:@3454.4]
  reg [63:0] _RAND_9;
  wire [63:0] tensorFile_4_1_rdata_4_data; // @[TensorLoad.scala 222:16:@3454.4]
  wire [9:0] tensorFile_4_1_rdata_4_addr; // @[TensorLoad.scala 222:16:@3454.4]
  wire [63:0] tensorFile_4_1__T_5324_data; // @[TensorLoad.scala 222:16:@3454.4]
  wire [9:0] tensorFile_4_1__T_5324_addr; // @[TensorLoad.scala 222:16:@3454.4]
  wire  tensorFile_4_1__T_5324_mask; // @[TensorLoad.scala 222:16:@3454.4]
  wire  tensorFile_4_1__T_5324_en; // @[TensorLoad.scala 222:16:@3454.4]
  reg [63:0] tensorFile_5_0 [0:1023]; // @[TensorLoad.scala 222:16:@3455.4]
  reg [63:0] _RAND_10;
  wire [63:0] tensorFile_5_0_rdata_5_data; // @[TensorLoad.scala 222:16:@3455.4]
  wire [9:0] tensorFile_5_0_rdata_5_addr; // @[TensorLoad.scala 222:16:@3455.4]
  wire [63:0] tensorFile_5_0__T_5411_data; // @[TensorLoad.scala 222:16:@3455.4]
  wire [9:0] tensorFile_5_0__T_5411_addr; // @[TensorLoad.scala 222:16:@3455.4]
  wire  tensorFile_5_0__T_5411_mask; // @[TensorLoad.scala 222:16:@3455.4]
  wire  tensorFile_5_0__T_5411_en; // @[TensorLoad.scala 222:16:@3455.4]
  reg [63:0] tensorFile_5_1 [0:1023]; // @[TensorLoad.scala 222:16:@3455.4]
  reg [63:0] _RAND_11;
  wire [63:0] tensorFile_5_1_rdata_5_data; // @[TensorLoad.scala 222:16:@3455.4]
  wire [9:0] tensorFile_5_1_rdata_5_addr; // @[TensorLoad.scala 222:16:@3455.4]
  wire [63:0] tensorFile_5_1__T_5411_data; // @[TensorLoad.scala 222:16:@3455.4]
  wire [9:0] tensorFile_5_1__T_5411_addr; // @[TensorLoad.scala 222:16:@3455.4]
  wire  tensorFile_5_1__T_5411_mask; // @[TensorLoad.scala 222:16:@3455.4]
  wire  tensorFile_5_1__T_5411_en; // @[TensorLoad.scala 222:16:@3455.4]
  reg [63:0] tensorFile_6_0 [0:1023]; // @[TensorLoad.scala 222:16:@3456.4]
  reg [63:0] _RAND_12;
  wire [63:0] tensorFile_6_0_rdata_6_data; // @[TensorLoad.scala 222:16:@3456.4]
  wire [9:0] tensorFile_6_0_rdata_6_addr; // @[TensorLoad.scala 222:16:@3456.4]
  wire [63:0] tensorFile_6_0__T_5498_data; // @[TensorLoad.scala 222:16:@3456.4]
  wire [9:0] tensorFile_6_0__T_5498_addr; // @[TensorLoad.scala 222:16:@3456.4]
  wire  tensorFile_6_0__T_5498_mask; // @[TensorLoad.scala 222:16:@3456.4]
  wire  tensorFile_6_0__T_5498_en; // @[TensorLoad.scala 222:16:@3456.4]
  reg [63:0] tensorFile_6_1 [0:1023]; // @[TensorLoad.scala 222:16:@3456.4]
  reg [63:0] _RAND_13;
  wire [63:0] tensorFile_6_1_rdata_6_data; // @[TensorLoad.scala 222:16:@3456.4]
  wire [9:0] tensorFile_6_1_rdata_6_addr; // @[TensorLoad.scala 222:16:@3456.4]
  wire [63:0] tensorFile_6_1__T_5498_data; // @[TensorLoad.scala 222:16:@3456.4]
  wire [9:0] tensorFile_6_1__T_5498_addr; // @[TensorLoad.scala 222:16:@3456.4]
  wire  tensorFile_6_1__T_5498_mask; // @[TensorLoad.scala 222:16:@3456.4]
  wire  tensorFile_6_1__T_5498_en; // @[TensorLoad.scala 222:16:@3456.4]
  reg [63:0] tensorFile_7_0 [0:1023]; // @[TensorLoad.scala 222:16:@3457.4]
  reg [63:0] _RAND_14;
  wire [63:0] tensorFile_7_0_rdata_7_data; // @[TensorLoad.scala 222:16:@3457.4]
  wire [9:0] tensorFile_7_0_rdata_7_addr; // @[TensorLoad.scala 222:16:@3457.4]
  wire [63:0] tensorFile_7_0__T_5585_data; // @[TensorLoad.scala 222:16:@3457.4]
  wire [9:0] tensorFile_7_0__T_5585_addr; // @[TensorLoad.scala 222:16:@3457.4]
  wire  tensorFile_7_0__T_5585_mask; // @[TensorLoad.scala 222:16:@3457.4]
  wire  tensorFile_7_0__T_5585_en; // @[TensorLoad.scala 222:16:@3457.4]
  reg [63:0] tensorFile_7_1 [0:1023]; // @[TensorLoad.scala 222:16:@3457.4]
  reg [63:0] _RAND_15;
  wire [63:0] tensorFile_7_1_rdata_7_data; // @[TensorLoad.scala 222:16:@3457.4]
  wire [9:0] tensorFile_7_1_rdata_7_addr; // @[TensorLoad.scala 222:16:@3457.4]
  wire [63:0] tensorFile_7_1__T_5585_data; // @[TensorLoad.scala 222:16:@3457.4]
  wire [9:0] tensorFile_7_1__T_5585_addr; // @[TensorLoad.scala 222:16:@3457.4]
  wire  tensorFile_7_1__T_5585_mask; // @[TensorLoad.scala 222:16:@3457.4]
  wire  tensorFile_7_1__T_5585_en; // @[TensorLoad.scala 222:16:@3457.4]
  reg [63:0] tensorFile_8_0 [0:1023]; // @[TensorLoad.scala 222:16:@3458.4]
  reg [63:0] _RAND_16;
  wire [63:0] tensorFile_8_0_rdata_8_data; // @[TensorLoad.scala 222:16:@3458.4]
  wire [9:0] tensorFile_8_0_rdata_8_addr; // @[TensorLoad.scala 222:16:@3458.4]
  wire [63:0] tensorFile_8_0__T_5672_data; // @[TensorLoad.scala 222:16:@3458.4]
  wire [9:0] tensorFile_8_0__T_5672_addr; // @[TensorLoad.scala 222:16:@3458.4]
  wire  tensorFile_8_0__T_5672_mask; // @[TensorLoad.scala 222:16:@3458.4]
  wire  tensorFile_8_0__T_5672_en; // @[TensorLoad.scala 222:16:@3458.4]
  reg [63:0] tensorFile_8_1 [0:1023]; // @[TensorLoad.scala 222:16:@3458.4]
  reg [63:0] _RAND_17;
  wire [63:0] tensorFile_8_1_rdata_8_data; // @[TensorLoad.scala 222:16:@3458.4]
  wire [9:0] tensorFile_8_1_rdata_8_addr; // @[TensorLoad.scala 222:16:@3458.4]
  wire [63:0] tensorFile_8_1__T_5672_data; // @[TensorLoad.scala 222:16:@3458.4]
  wire [9:0] tensorFile_8_1__T_5672_addr; // @[TensorLoad.scala 222:16:@3458.4]
  wire  tensorFile_8_1__T_5672_mask; // @[TensorLoad.scala 222:16:@3458.4]
  wire  tensorFile_8_1__T_5672_en; // @[TensorLoad.scala 222:16:@3458.4]
  reg [63:0] tensorFile_9_0 [0:1023]; // @[TensorLoad.scala 222:16:@3459.4]
  reg [63:0] _RAND_18;
  wire [63:0] tensorFile_9_0_rdata_9_data; // @[TensorLoad.scala 222:16:@3459.4]
  wire [9:0] tensorFile_9_0_rdata_9_addr; // @[TensorLoad.scala 222:16:@3459.4]
  wire [63:0] tensorFile_9_0__T_5759_data; // @[TensorLoad.scala 222:16:@3459.4]
  wire [9:0] tensorFile_9_0__T_5759_addr; // @[TensorLoad.scala 222:16:@3459.4]
  wire  tensorFile_9_0__T_5759_mask; // @[TensorLoad.scala 222:16:@3459.4]
  wire  tensorFile_9_0__T_5759_en; // @[TensorLoad.scala 222:16:@3459.4]
  reg [63:0] tensorFile_9_1 [0:1023]; // @[TensorLoad.scala 222:16:@3459.4]
  reg [63:0] _RAND_19;
  wire [63:0] tensorFile_9_1_rdata_9_data; // @[TensorLoad.scala 222:16:@3459.4]
  wire [9:0] tensorFile_9_1_rdata_9_addr; // @[TensorLoad.scala 222:16:@3459.4]
  wire [63:0] tensorFile_9_1__T_5759_data; // @[TensorLoad.scala 222:16:@3459.4]
  wire [9:0] tensorFile_9_1__T_5759_addr; // @[TensorLoad.scala 222:16:@3459.4]
  wire  tensorFile_9_1__T_5759_mask; // @[TensorLoad.scala 222:16:@3459.4]
  wire  tensorFile_9_1__T_5759_en; // @[TensorLoad.scala 222:16:@3459.4]
  reg [63:0] tensorFile_10_0 [0:1023]; // @[TensorLoad.scala 222:16:@3460.4]
  reg [63:0] _RAND_20;
  wire [63:0] tensorFile_10_0_rdata_10_data; // @[TensorLoad.scala 222:16:@3460.4]
  wire [9:0] tensorFile_10_0_rdata_10_addr; // @[TensorLoad.scala 222:16:@3460.4]
  wire [63:0] tensorFile_10_0__T_5846_data; // @[TensorLoad.scala 222:16:@3460.4]
  wire [9:0] tensorFile_10_0__T_5846_addr; // @[TensorLoad.scala 222:16:@3460.4]
  wire  tensorFile_10_0__T_5846_mask; // @[TensorLoad.scala 222:16:@3460.4]
  wire  tensorFile_10_0__T_5846_en; // @[TensorLoad.scala 222:16:@3460.4]
  reg [63:0] tensorFile_10_1 [0:1023]; // @[TensorLoad.scala 222:16:@3460.4]
  reg [63:0] _RAND_21;
  wire [63:0] tensorFile_10_1_rdata_10_data; // @[TensorLoad.scala 222:16:@3460.4]
  wire [9:0] tensorFile_10_1_rdata_10_addr; // @[TensorLoad.scala 222:16:@3460.4]
  wire [63:0] tensorFile_10_1__T_5846_data; // @[TensorLoad.scala 222:16:@3460.4]
  wire [9:0] tensorFile_10_1__T_5846_addr; // @[TensorLoad.scala 222:16:@3460.4]
  wire  tensorFile_10_1__T_5846_mask; // @[TensorLoad.scala 222:16:@3460.4]
  wire  tensorFile_10_1__T_5846_en; // @[TensorLoad.scala 222:16:@3460.4]
  reg [63:0] tensorFile_11_0 [0:1023]; // @[TensorLoad.scala 222:16:@3461.4]
  reg [63:0] _RAND_22;
  wire [63:0] tensorFile_11_0_rdata_11_data; // @[TensorLoad.scala 222:16:@3461.4]
  wire [9:0] tensorFile_11_0_rdata_11_addr; // @[TensorLoad.scala 222:16:@3461.4]
  wire [63:0] tensorFile_11_0__T_5933_data; // @[TensorLoad.scala 222:16:@3461.4]
  wire [9:0] tensorFile_11_0__T_5933_addr; // @[TensorLoad.scala 222:16:@3461.4]
  wire  tensorFile_11_0__T_5933_mask; // @[TensorLoad.scala 222:16:@3461.4]
  wire  tensorFile_11_0__T_5933_en; // @[TensorLoad.scala 222:16:@3461.4]
  reg [63:0] tensorFile_11_1 [0:1023]; // @[TensorLoad.scala 222:16:@3461.4]
  reg [63:0] _RAND_23;
  wire [63:0] tensorFile_11_1_rdata_11_data; // @[TensorLoad.scala 222:16:@3461.4]
  wire [9:0] tensorFile_11_1_rdata_11_addr; // @[TensorLoad.scala 222:16:@3461.4]
  wire [63:0] tensorFile_11_1__T_5933_data; // @[TensorLoad.scala 222:16:@3461.4]
  wire [9:0] tensorFile_11_1__T_5933_addr; // @[TensorLoad.scala 222:16:@3461.4]
  wire  tensorFile_11_1__T_5933_mask; // @[TensorLoad.scala 222:16:@3461.4]
  wire  tensorFile_11_1__T_5933_en; // @[TensorLoad.scala 222:16:@3461.4]
  reg [63:0] tensorFile_12_0 [0:1023]; // @[TensorLoad.scala 222:16:@3462.4]
  reg [63:0] _RAND_24;
  wire [63:0] tensorFile_12_0_rdata_12_data; // @[TensorLoad.scala 222:16:@3462.4]
  wire [9:0] tensorFile_12_0_rdata_12_addr; // @[TensorLoad.scala 222:16:@3462.4]
  wire [63:0] tensorFile_12_0__T_6020_data; // @[TensorLoad.scala 222:16:@3462.4]
  wire [9:0] tensorFile_12_0__T_6020_addr; // @[TensorLoad.scala 222:16:@3462.4]
  wire  tensorFile_12_0__T_6020_mask; // @[TensorLoad.scala 222:16:@3462.4]
  wire  tensorFile_12_0__T_6020_en; // @[TensorLoad.scala 222:16:@3462.4]
  reg [63:0] tensorFile_12_1 [0:1023]; // @[TensorLoad.scala 222:16:@3462.4]
  reg [63:0] _RAND_25;
  wire [63:0] tensorFile_12_1_rdata_12_data; // @[TensorLoad.scala 222:16:@3462.4]
  wire [9:0] tensorFile_12_1_rdata_12_addr; // @[TensorLoad.scala 222:16:@3462.4]
  wire [63:0] tensorFile_12_1__T_6020_data; // @[TensorLoad.scala 222:16:@3462.4]
  wire [9:0] tensorFile_12_1__T_6020_addr; // @[TensorLoad.scala 222:16:@3462.4]
  wire  tensorFile_12_1__T_6020_mask; // @[TensorLoad.scala 222:16:@3462.4]
  wire  tensorFile_12_1__T_6020_en; // @[TensorLoad.scala 222:16:@3462.4]
  reg [63:0] tensorFile_13_0 [0:1023]; // @[TensorLoad.scala 222:16:@3463.4]
  reg [63:0] _RAND_26;
  wire [63:0] tensorFile_13_0_rdata_13_data; // @[TensorLoad.scala 222:16:@3463.4]
  wire [9:0] tensorFile_13_0_rdata_13_addr; // @[TensorLoad.scala 222:16:@3463.4]
  wire [63:0] tensorFile_13_0__T_6107_data; // @[TensorLoad.scala 222:16:@3463.4]
  wire [9:0] tensorFile_13_0__T_6107_addr; // @[TensorLoad.scala 222:16:@3463.4]
  wire  tensorFile_13_0__T_6107_mask; // @[TensorLoad.scala 222:16:@3463.4]
  wire  tensorFile_13_0__T_6107_en; // @[TensorLoad.scala 222:16:@3463.4]
  reg [63:0] tensorFile_13_1 [0:1023]; // @[TensorLoad.scala 222:16:@3463.4]
  reg [63:0] _RAND_27;
  wire [63:0] tensorFile_13_1_rdata_13_data; // @[TensorLoad.scala 222:16:@3463.4]
  wire [9:0] tensorFile_13_1_rdata_13_addr; // @[TensorLoad.scala 222:16:@3463.4]
  wire [63:0] tensorFile_13_1__T_6107_data; // @[TensorLoad.scala 222:16:@3463.4]
  wire [9:0] tensorFile_13_1__T_6107_addr; // @[TensorLoad.scala 222:16:@3463.4]
  wire  tensorFile_13_1__T_6107_mask; // @[TensorLoad.scala 222:16:@3463.4]
  wire  tensorFile_13_1__T_6107_en; // @[TensorLoad.scala 222:16:@3463.4]
  reg [63:0] tensorFile_14_0 [0:1023]; // @[TensorLoad.scala 222:16:@3464.4]
  reg [63:0] _RAND_28;
  wire [63:0] tensorFile_14_0_rdata_14_data; // @[TensorLoad.scala 222:16:@3464.4]
  wire [9:0] tensorFile_14_0_rdata_14_addr; // @[TensorLoad.scala 222:16:@3464.4]
  wire [63:0] tensorFile_14_0__T_6194_data; // @[TensorLoad.scala 222:16:@3464.4]
  wire [9:0] tensorFile_14_0__T_6194_addr; // @[TensorLoad.scala 222:16:@3464.4]
  wire  tensorFile_14_0__T_6194_mask; // @[TensorLoad.scala 222:16:@3464.4]
  wire  tensorFile_14_0__T_6194_en; // @[TensorLoad.scala 222:16:@3464.4]
  reg [63:0] tensorFile_14_1 [0:1023]; // @[TensorLoad.scala 222:16:@3464.4]
  reg [63:0] _RAND_29;
  wire [63:0] tensorFile_14_1_rdata_14_data; // @[TensorLoad.scala 222:16:@3464.4]
  wire [9:0] tensorFile_14_1_rdata_14_addr; // @[TensorLoad.scala 222:16:@3464.4]
  wire [63:0] tensorFile_14_1__T_6194_data; // @[TensorLoad.scala 222:16:@3464.4]
  wire [9:0] tensorFile_14_1__T_6194_addr; // @[TensorLoad.scala 222:16:@3464.4]
  wire  tensorFile_14_1__T_6194_mask; // @[TensorLoad.scala 222:16:@3464.4]
  wire  tensorFile_14_1__T_6194_en; // @[TensorLoad.scala 222:16:@3464.4]
  reg [63:0] tensorFile_15_0 [0:1023]; // @[TensorLoad.scala 222:16:@3465.4]
  reg [63:0] _RAND_30;
  wire [63:0] tensorFile_15_0_rdata_15_data; // @[TensorLoad.scala 222:16:@3465.4]
  wire [9:0] tensorFile_15_0_rdata_15_addr; // @[TensorLoad.scala 222:16:@3465.4]
  wire [63:0] tensorFile_15_0__T_6281_data; // @[TensorLoad.scala 222:16:@3465.4]
  wire [9:0] tensorFile_15_0__T_6281_addr; // @[TensorLoad.scala 222:16:@3465.4]
  wire  tensorFile_15_0__T_6281_mask; // @[TensorLoad.scala 222:16:@3465.4]
  wire  tensorFile_15_0__T_6281_en; // @[TensorLoad.scala 222:16:@3465.4]
  reg [63:0] tensorFile_15_1 [0:1023]; // @[TensorLoad.scala 222:16:@3465.4]
  reg [63:0] _RAND_31;
  wire [63:0] tensorFile_15_1_rdata_15_data; // @[TensorLoad.scala 222:16:@3465.4]
  wire [9:0] tensorFile_15_1_rdata_15_addr; // @[TensorLoad.scala 222:16:@3465.4]
  wire [63:0] tensorFile_15_1__T_6281_data; // @[TensorLoad.scala 222:16:@3465.4]
  wire [9:0] tensorFile_15_1__T_6281_addr; // @[TensorLoad.scala 222:16:@3465.4]
  wire  tensorFile_15_1__T_6281_mask; // @[TensorLoad.scala 222:16:@3465.4]
  wire  tensorFile_15_1__T_6281_en; // @[TensorLoad.scala 222:16:@3465.4]
  wire [15:0] dec_sram_offset; // @[TensorLoad.scala 51:29:@3147.4]
  wire [15:0] dec_xsize; // @[TensorLoad.scala 51:29:@3155.4]
  wire [3:0] dec_ypad_0; // @[TensorLoad.scala 51:29:@3159.4]
  wire [3:0] dec_ypad_1; // @[TensorLoad.scala 51:29:@3161.4]
  wire [3:0] dec_xpad_0; // @[TensorLoad.scala 51:29:@3163.4]
  wire [3:0] dec_xpad_1; // @[TensorLoad.scala 51:29:@3165.4]
  reg  dataCtrlDone; // @[TensorLoad.scala 54:29:@3170.4]
  reg [31:0] _RAND_32;
  reg  tag; // @[TensorLoad.scala 60:16:@3183.4]
  reg [31:0] _RAND_33;
  reg [3:0] set; // @[TensorLoad.scala 61:16:@3184.4]
  reg [31:0] _RAND_34;
  reg [2:0] state; // @[TensorLoad.scala 65:22:@3185.4]
  reg [31:0] _RAND_35;
  wire  _T_4394; // @[Conditional.scala 37:30:@3186.4]
  wire  _T_4396; // @[TensorLoad.scala 71:25:@3189.8]
  wire  _T_4398; // @[TensorLoad.scala 73:31:@3194.10]
  wire [2:0] _GEN_0; // @[TensorLoad.scala 73:40:@3195.10]
  wire [2:0] _GEN_1; // @[TensorLoad.scala 71:34:@3190.8]
  wire [2:0] _GEN_2; // @[TensorLoad.scala 70:22:@3188.6]
  wire  _T_4399; // @[Conditional.scala 37:30:@3204.6]
  wire [2:0] _GEN_4; // @[TensorLoad.scala 81:31:@3206.8]
  wire  _T_4402; // @[Conditional.scala 37:30:@3217.8]
  wire [2:0] _GEN_5; // @[TensorLoad.scala 90:31:@3219.10]
  wire  _T_4403; // @[Conditional.scala 37:30:@3224.10]
  wire [2:0] _GEN_6; // @[TensorLoad.scala 95:33:@3226.12]
  wire  _T_4404; // @[Conditional.scala 37:30:@3231.12]
  wire  _T_4406; // @[TensorLoad.scala 102:27:@3235.18]
  wire  _T_4408; // @[TensorLoad.scala 104:33:@3240.20]
  wire [2:0] _GEN_7; // @[TensorLoad.scala 104:42:@3241.20]
  wire [2:0] _GEN_8; // @[TensorLoad.scala 102:36:@3236.18]
  wire [2:0] _GEN_10; // @[TensorLoad.scala 110:36:@3251.20]
  wire [2:0] _GEN_11; // @[TensorLoad.scala 117:39:@3264.20]
  wire [2:0] _GEN_12; // @[TensorLoad.scala 109:40:@3249.18]
  wire [2:0] _GEN_13; // @[TensorLoad.scala 101:32:@3234.16]
  wire [2:0] _GEN_14; // @[TensorLoad.scala 100:34:@3233.14]
  wire  _T_4413; // @[Conditional.scala 37:30:@3270.14]
  wire [2:0] _GEN_17; // @[TensorLoad.scala 124:28:@3273.18]
  wire [2:0] _GEN_18; // @[TensorLoad.scala 123:31:@3272.16]
  wire  _T_4418; // @[Conditional.scala 37:30:@3294.16]
  wire  _T_4419; // @[TensorLoad.scala 140:30:@3296.18]
  wire [2:0] _GEN_19; // @[TensorLoad.scala 140:47:@3297.18]
  wire [2:0] _GEN_20; // @[Conditional.scala 39:67:@3295.16]
  wire [2:0] _GEN_21; // @[Conditional.scala 39:67:@3271.14]
  wire [2:0] _GEN_22; // @[Conditional.scala 39:67:@3232.12]
  wire [2:0] _GEN_23; // @[Conditional.scala 39:67:@3225.10]
  wire [2:0] _GEN_24; // @[Conditional.scala 39:67:@3218.8]
  wire [2:0] _GEN_25; // @[Conditional.scala 39:67:@3205.6]
  wire [2:0] _GEN_26; // @[Conditional.scala 40:58:@3187.4]
  wire  _T_4420; // @[TensorLoad.scala 147:30:@3301.4]
  wire  _T_4421; // @[TensorLoad.scala 147:40:@3302.4]
  wire  _T_4423; // @[Decoupled.scala 37:37:@3308.4]
  wire  _T_4428; // @[TensorLoad.scala 156:36:@3318.6]
  wire  _GEN_27; // @[TensorLoad.scala 156:57:@3319.6]
  wire  _GEN_28; // @[TensorLoad.scala 154:25:@3313.4]
  wire  _T_4433; // @[TensorLoad.scala 161:44:@3324.4]
  wire  _T_4440; // @[TensorLoad.scala 164:61:@3330.4]
  wire  _T_4441; // @[TensorLoad.scala 164:48:@3331.4]
  wire  _T_4442; // @[TensorLoad.scala 165:14:@3332.4]
  wire  _T_4443; // @[TensorLoad.scala 165:25:@3333.4]
  wire  _T_4444; // @[TensorLoad.scala 165:45:@3334.4]
  wire  _T_4445; // @[TensorLoad.scala 164:70:@3335.4]
  wire  _T_4451; // @[TensorLoad.scala 169:14:@3341.4]
  wire  _T_4452; // @[TensorLoad.scala 169:25:@3342.4]
  wire  _T_4453; // @[TensorLoad.scala 168:35:@3343.4]
  wire  _T_4455; // @[TensorLoad.scala 170:32:@3345.4]
  wire  _T_4456; // @[TensorLoad.scala 170:30:@3346.4]
  wire  _T_4457; // @[TensorLoad.scala 170:46:@3347.4]
  wire  _T_4460; // @[TensorLoad.scala 170:67:@3349.4]
  wire  _T_4461; // @[TensorLoad.scala 169:46:@3350.4]
  wire  _T_4465; // @[TensorLoad.scala 171:45:@3354.4]
  wire  _T_4466; // @[TensorLoad.scala 170:89:@3355.4]
  wire  _T_4471; // @[TensorLoad.scala 173:44:@3360.4]
  wire  _T_4472; // @[TensorLoad.scala 174:28:@3361.4]
  wire  _T_4473; // @[TensorLoad.scala 174:46:@3362.4]
  wire  _T_4476; // @[TensorLoad.scala 174:67:@3364.4]
  wire  _T_4477; // @[TensorLoad.scala 174:25:@3365.4]
  wire  _T_4479; // @[TensorLoad.scala 182:32:@3372.4]
  wire  _T_4482; // @[TensorLoad.scala 190:11:@3379.4]
  wire  _T_4483; // @[TensorLoad.scala 189:36:@3380.4]
  wire  _T_4485; // @[TensorLoad.scala 190:22:@3382.4]
  wire  _T_4486; // @[TensorLoad.scala 192:11:@3383.4]
  wire  isZeroPad; // @[TensorLoad.scala 191:22:@3384.4]
  wire  _T_4489; // @[TensorLoad.scala 194:24:@3387.4]
  wire  _T_4492; // @[TensorLoad.scala 194:46:@3389.4]
  wire  _T_4495; // @[TensorLoad.scala 196:36:@3395.6]
  wire [1:0] _T_4497; // @[TensorLoad.scala 197:16:@3397.8]
  wire  _T_4498; // @[TensorLoad.scala 197:16:@3398.8]
  wire  _GEN_29; // @[TensorLoad.scala 196:50:@3396.6]
  wire  _T_4500; // @[TensorLoad.scala 200:24:@3402.4]
  wire  _T_4502; // @[TensorLoad.scala 200:48:@3403.4]
  wire  _T_4505; // @[TensorLoad.scala 200:76:@3405.4]
  wire  _T_4506; // @[TensorLoad.scala 200:40:@3406.4]
  wire  _T_4512; // @[TensorLoad.scala 202:51:@3414.6]
  wire [4:0] _T_4514; // @[TensorLoad.scala 203:16:@3416.8]
  wire [3:0] _T_4515; // @[TensorLoad.scala 203:16:@3417.8]
  wire [3:0] _GEN_31; // @[TensorLoad.scala 202:86:@3415.6]
  reg [9:0] waddr_cur; // @[TensorLoad.scala 206:22:@3420.4]
  reg [31:0] _RAND_36;
  reg [9:0] waddr_nxt; // @[TensorLoad.scala 207:22:@3421.4]
  reg [31:0] _RAND_37;
  wire  _T_4523; // @[TensorLoad.scala 212:5:@3431.6]
  wire  _T_4526; // @[TensorLoad.scala 213:5:@3433.6]
  wire [10:0] _T_4528; // @[TensorLoad.scala 215:28:@3435.8]
  wire [9:0] _T_4529; // @[TensorLoad.scala 215:28:@3436.8]
  wire  _T_4531; // @[TensorLoad.scala 216:33:@3441.8]
  wire [15:0] _GEN_426; // @[TensorLoad.scala 217:28:@3443.10]
  wire [16:0] _T_4532; // @[TensorLoad.scala 217:28:@3443.10]
  wire [15:0] _T_4533; // @[TensorLoad.scala 217:28:@3444.10]
  wire [15:0] _GEN_33; // @[TensorLoad.scala 216:59:@3442.8]
  wire [15:0] _GEN_34; // @[TensorLoad.scala 216:59:@3442.8]
  wire [15:0] _GEN_35; // @[TensorLoad.scala 214:3:@3434.6]
  wire [15:0] _GEN_36; // @[TensorLoad.scala 214:3:@3434.6]
  wire [15:0] _GEN_37; // @[TensorLoad.scala 208:25:@3423.4]
  wire [15:0] _GEN_38; // @[TensorLoad.scala 208:25:@3423.4]
  wire  wmask_0_0; // @[TensorLoad.scala 235:26:@3501.4]
  wire [63:0] wdata_0_0; // @[TensorLoad.scala 236:25:@3503.4]
  wire  _T_4947; // @[TensorLoad.scala 242:51:@3534.4]
  wire  _T_4948; // @[TensorLoad.scala 242:45:@3535.4]
  wire  _T_5034; // @[TensorLoad.scala 242:51:@3585.4]
  wire  _T_5035; // @[TensorLoad.scala 242:45:@3586.4]
  wire  _T_5121; // @[TensorLoad.scala 242:51:@3636.4]
  wire  _T_5122; // @[TensorLoad.scala 242:45:@3637.4]
  wire  _T_5208; // @[TensorLoad.scala 242:51:@3687.4]
  wire  _T_5209; // @[TensorLoad.scala 242:45:@3688.4]
  wire  _T_5295; // @[TensorLoad.scala 242:51:@3738.4]
  wire  _T_5296; // @[TensorLoad.scala 242:45:@3739.4]
  wire  _T_5382; // @[TensorLoad.scala 242:51:@3789.4]
  wire  _T_5383; // @[TensorLoad.scala 242:45:@3790.4]
  wire  _T_5469; // @[TensorLoad.scala 242:51:@3840.4]
  wire  _T_5470; // @[TensorLoad.scala 242:45:@3841.4]
  wire  _T_5556; // @[TensorLoad.scala 242:51:@3891.4]
  wire  _T_5557; // @[TensorLoad.scala 242:45:@3892.4]
  wire  _T_5643; // @[TensorLoad.scala 242:51:@3942.4]
  wire  _T_5644; // @[TensorLoad.scala 242:45:@3943.4]
  wire  _T_5730; // @[TensorLoad.scala 242:51:@3993.4]
  wire  _T_5731; // @[TensorLoad.scala 242:45:@3994.4]
  wire  _T_5817; // @[TensorLoad.scala 242:51:@4044.4]
  wire  _T_5818; // @[TensorLoad.scala 242:45:@4045.4]
  wire  _T_5904; // @[TensorLoad.scala 242:51:@4095.4]
  wire  _T_5905; // @[TensorLoad.scala 242:45:@4096.4]
  wire  _T_5991; // @[TensorLoad.scala 242:51:@4146.4]
  wire  _T_5992; // @[TensorLoad.scala 242:45:@4147.4]
  wire  _T_6078; // @[TensorLoad.scala 242:51:@4197.4]
  wire  _T_6079; // @[TensorLoad.scala 242:45:@4198.4]
  wire  _T_6165; // @[TensorLoad.scala 242:51:@4248.4]
  wire  _T_6166; // @[TensorLoad.scala 242:45:@4249.4]
  reg  rvalid; // @[TensorLoad.scala 252:23:@4317.4]
  reg [31:0] _RAND_38;
  wire  _GEN_216; // @[TensorLoad.scala 256:26:@4322.4]
  wire [127:0] _T_6482; // @[TensorLoad.scala 259:38:@4448.4]
  wire [127:0] _T_6624; // @[TensorLoad.scala 259:38:@4500.4]
  wire [127:0] _T_6766; // @[TensorLoad.scala 259:38:@4552.4]
  wire [127:0] _T_6908; // @[TensorLoad.scala 259:38:@4604.4]
  wire [127:0] _T_7050; // @[TensorLoad.scala 259:38:@4656.4]
  wire [127:0] _T_7192; // @[TensorLoad.scala 259:38:@4708.4]
  wire [127:0] _T_7334; // @[TensorLoad.scala 259:38:@4760.4]
  wire [127:0] _T_7476; // @[TensorLoad.scala 259:38:@4812.4]
  wire [127:0] _T_7618; // @[TensorLoad.scala 259:38:@4864.4]
  wire [127:0] _T_7760; // @[TensorLoad.scala 259:38:@4916.4]
  wire [127:0] _T_7902; // @[TensorLoad.scala 259:38:@4968.4]
  wire [127:0] _T_8044; // @[TensorLoad.scala 259:38:@5020.4]
  wire [127:0] _T_8186; // @[TensorLoad.scala 259:38:@5072.4]
  wire [127:0] _T_8328; // @[TensorLoad.scala 259:38:@5124.4]
  wire [127:0] _T_8470; // @[TensorLoad.scala 259:38:@5176.4]
  wire [127:0] _T_8612; // @[TensorLoad.scala 259:38:@5228.4]
  wire  _T_8760; // @[TensorLoad.scala 263:96:@5284.4]
  wire  done_no_pad; // @[TensorLoad.scala 263:83:@5285.4]
  wire  done_x_pad; // @[TensorLoad.scala 264:72:@5290.4]
  wire  _T_8767; // @[TensorLoad.scala 265:37:@5292.4]
  wire  done_y_pad; // @[TensorLoad.scala 265:52:@5293.4]
  wire  _T_8768; // @[TensorLoad.scala 266:26:@5294.4]
  reg [9:0] tensorFile_0_0_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_39;
  reg [9:0] tensorFile_0_1_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_40;
  reg [9:0] tensorFile_1_0_rdata_1_addr_pipe_0;
  reg [31:0] _RAND_41;
  reg [9:0] tensorFile_1_1_rdata_1_addr_pipe_0;
  reg [31:0] _RAND_42;
  reg [9:0] tensorFile_2_0_rdata_2_addr_pipe_0;
  reg [31:0] _RAND_43;
  reg [9:0] tensorFile_2_1_rdata_2_addr_pipe_0;
  reg [31:0] _RAND_44;
  reg [9:0] tensorFile_3_0_rdata_3_addr_pipe_0;
  reg [31:0] _RAND_45;
  reg [9:0] tensorFile_3_1_rdata_3_addr_pipe_0;
  reg [31:0] _RAND_46;
  reg [9:0] tensorFile_4_0_rdata_4_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [9:0] tensorFile_4_1_rdata_4_addr_pipe_0;
  reg [31:0] _RAND_48;
  reg [9:0] tensorFile_5_0_rdata_5_addr_pipe_0;
  reg [31:0] _RAND_49;
  reg [9:0] tensorFile_5_1_rdata_5_addr_pipe_0;
  reg [31:0] _RAND_50;
  reg [9:0] tensorFile_6_0_rdata_6_addr_pipe_0;
  reg [31:0] _RAND_51;
  reg [9:0] tensorFile_6_1_rdata_6_addr_pipe_0;
  reg [31:0] _RAND_52;
  reg [9:0] tensorFile_7_0_rdata_7_addr_pipe_0;
  reg [31:0] _RAND_53;
  reg [9:0] tensorFile_7_1_rdata_7_addr_pipe_0;
  reg [31:0] _RAND_54;
  reg [9:0] tensorFile_8_0_rdata_8_addr_pipe_0;
  reg [31:0] _RAND_55;
  reg [9:0] tensorFile_8_1_rdata_8_addr_pipe_0;
  reg [31:0] _RAND_56;
  reg [9:0] tensorFile_9_0_rdata_9_addr_pipe_0;
  reg [31:0] _RAND_57;
  reg [9:0] tensorFile_9_1_rdata_9_addr_pipe_0;
  reg [31:0] _RAND_58;
  reg [9:0] tensorFile_10_0_rdata_10_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [9:0] tensorFile_10_1_rdata_10_addr_pipe_0;
  reg [31:0] _RAND_60;
  reg [9:0] tensorFile_11_0_rdata_11_addr_pipe_0;
  reg [31:0] _RAND_61;
  reg [9:0] tensorFile_11_1_rdata_11_addr_pipe_0;
  reg [31:0] _RAND_62;
  reg [9:0] tensorFile_12_0_rdata_12_addr_pipe_0;
  reg [31:0] _RAND_63;
  reg [9:0] tensorFile_12_1_rdata_12_addr_pipe_0;
  reg [31:0] _RAND_64;
  reg [9:0] tensorFile_13_0_rdata_13_addr_pipe_0;
  reg [31:0] _RAND_65;
  reg [9:0] tensorFile_13_1_rdata_13_addr_pipe_0;
  reg [31:0] _RAND_66;
  reg [9:0] tensorFile_14_0_rdata_14_addr_pipe_0;
  reg [31:0] _RAND_67;
  reg [9:0] tensorFile_14_1_rdata_14_addr_pipe_0;
  reg [31:0] _RAND_68;
  reg [9:0] tensorFile_15_0_rdata_15_addr_pipe_0;
  reg [31:0] _RAND_69;
  reg [9:0] tensorFile_15_1_rdata_15_addr_pipe_0;
  reg [31:0] _RAND_70;
  TensorDataCtrl_1 dataCtrl ( // @[TensorLoad.scala 52:24:@3167.4]
    .clock(dataCtrl_clock),
    .io_start(dataCtrl_io_start),
    .io_done(dataCtrl_io_done),
    .io_inst(dataCtrl_io_inst),
    .io_baddr(dataCtrl_io_baddr),
    .io_xinit(dataCtrl_io_xinit),
    .io_xupdate(dataCtrl_io_xupdate),
    .io_yupdate(dataCtrl_io_yupdate),
    .io_stride(dataCtrl_io_stride),
    .io_split(dataCtrl_io_split),
    .io_addr(dataCtrl_io_addr),
    .io_len(dataCtrl_io_len)
  );
  TensorPadCtrl_4 yPadCtrl0 ( // @[TensorLoad.scala 55:25:@3171.4]
    .clock(yPadCtrl0_clock),
    .reset(yPadCtrl0_reset),
    .io_start(yPadCtrl0_io_start),
    .io_done(yPadCtrl0_io_done),
    .io_inst(yPadCtrl0_io_inst)
  );
  TensorPadCtrl_5 yPadCtrl1 ( // @[TensorLoad.scala 56:25:@3174.4]
    .clock(yPadCtrl1_clock),
    .reset(yPadCtrl1_reset),
    .io_start(yPadCtrl1_io_start),
    .io_done(yPadCtrl1_io_done),
    .io_inst(yPadCtrl1_io_inst)
  );
  TensorPadCtrl_6 xPadCtrl0 ( // @[TensorLoad.scala 57:25:@3177.4]
    .clock(xPadCtrl0_clock),
    .reset(xPadCtrl0_reset),
    .io_start(xPadCtrl0_io_start),
    .io_done(xPadCtrl0_io_done),
    .io_inst(xPadCtrl0_io_inst)
  );
  TensorPadCtrl_7 xPadCtrl1 ( // @[TensorLoad.scala 58:25:@3180.4]
    .clock(xPadCtrl1_clock),
    .reset(xPadCtrl1_reset),
    .io_start(xPadCtrl1_io_start),
    .io_done(xPadCtrl1_io_done),
    .io_inst(xPadCtrl1_io_inst)
  );
  assign tensorFile_0_0_rdata_0_addr = tensorFile_0_0_rdata_0_addr_pipe_0;
  assign tensorFile_0_0_rdata_0_data = tensorFile_0_0[tensorFile_0_0_rdata_0_addr]; // @[TensorLoad.scala 222:16:@3450.4]
  assign tensorFile_0_0__T_4976_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_0_0__T_4976_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_0_0__T_4976_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_0_0__T_4976_en = _T_4420 ? 1'h0 : _T_4948;
  assign tensorFile_0_1_rdata_0_addr = tensorFile_0_1_rdata_0_addr_pipe_0;
  assign tensorFile_0_1_rdata_0_data = tensorFile_0_1[tensorFile_0_1_rdata_0_addr]; // @[TensorLoad.scala 222:16:@3450.4]
  assign tensorFile_0_1__T_4976_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_0_1__T_4976_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_0_1__T_4976_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_0_1__T_4976_en = _T_4420 ? 1'h0 : _T_4948;
  assign tensorFile_1_0_rdata_1_addr = tensorFile_1_0_rdata_1_addr_pipe_0;
  assign tensorFile_1_0_rdata_1_data = tensorFile_1_0[tensorFile_1_0_rdata_1_addr]; // @[TensorLoad.scala 222:16:@3451.4]
  assign tensorFile_1_0__T_5063_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_1_0__T_5063_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_1_0__T_5063_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_1_0__T_5063_en = _T_4420 ? 1'h0 : _T_5035;
  assign tensorFile_1_1_rdata_1_addr = tensorFile_1_1_rdata_1_addr_pipe_0;
  assign tensorFile_1_1_rdata_1_data = tensorFile_1_1[tensorFile_1_1_rdata_1_addr]; // @[TensorLoad.scala 222:16:@3451.4]
  assign tensorFile_1_1__T_5063_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_1_1__T_5063_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_1_1__T_5063_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_1_1__T_5063_en = _T_4420 ? 1'h0 : _T_5035;
  assign tensorFile_2_0_rdata_2_addr = tensorFile_2_0_rdata_2_addr_pipe_0;
  assign tensorFile_2_0_rdata_2_data = tensorFile_2_0[tensorFile_2_0_rdata_2_addr]; // @[TensorLoad.scala 222:16:@3452.4]
  assign tensorFile_2_0__T_5150_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_2_0__T_5150_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_2_0__T_5150_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_2_0__T_5150_en = _T_4420 ? 1'h0 : _T_5122;
  assign tensorFile_2_1_rdata_2_addr = tensorFile_2_1_rdata_2_addr_pipe_0;
  assign tensorFile_2_1_rdata_2_data = tensorFile_2_1[tensorFile_2_1_rdata_2_addr]; // @[TensorLoad.scala 222:16:@3452.4]
  assign tensorFile_2_1__T_5150_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_2_1__T_5150_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_2_1__T_5150_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_2_1__T_5150_en = _T_4420 ? 1'h0 : _T_5122;
  assign tensorFile_3_0_rdata_3_addr = tensorFile_3_0_rdata_3_addr_pipe_0;
  assign tensorFile_3_0_rdata_3_data = tensorFile_3_0[tensorFile_3_0_rdata_3_addr]; // @[TensorLoad.scala 222:16:@3453.4]
  assign tensorFile_3_0__T_5237_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_3_0__T_5237_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_3_0__T_5237_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_3_0__T_5237_en = _T_4420 ? 1'h0 : _T_5209;
  assign tensorFile_3_1_rdata_3_addr = tensorFile_3_1_rdata_3_addr_pipe_0;
  assign tensorFile_3_1_rdata_3_data = tensorFile_3_1[tensorFile_3_1_rdata_3_addr]; // @[TensorLoad.scala 222:16:@3453.4]
  assign tensorFile_3_1__T_5237_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_3_1__T_5237_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_3_1__T_5237_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_3_1__T_5237_en = _T_4420 ? 1'h0 : _T_5209;
  assign tensorFile_4_0_rdata_4_addr = tensorFile_4_0_rdata_4_addr_pipe_0;
  assign tensorFile_4_0_rdata_4_data = tensorFile_4_0[tensorFile_4_0_rdata_4_addr]; // @[TensorLoad.scala 222:16:@3454.4]
  assign tensorFile_4_0__T_5324_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_4_0__T_5324_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_4_0__T_5324_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_4_0__T_5324_en = _T_4420 ? 1'h0 : _T_5296;
  assign tensorFile_4_1_rdata_4_addr = tensorFile_4_1_rdata_4_addr_pipe_0;
  assign tensorFile_4_1_rdata_4_data = tensorFile_4_1[tensorFile_4_1_rdata_4_addr]; // @[TensorLoad.scala 222:16:@3454.4]
  assign tensorFile_4_1__T_5324_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_4_1__T_5324_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_4_1__T_5324_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_4_1__T_5324_en = _T_4420 ? 1'h0 : _T_5296;
  assign tensorFile_5_0_rdata_5_addr = tensorFile_5_0_rdata_5_addr_pipe_0;
  assign tensorFile_5_0_rdata_5_data = tensorFile_5_0[tensorFile_5_0_rdata_5_addr]; // @[TensorLoad.scala 222:16:@3455.4]
  assign tensorFile_5_0__T_5411_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_5_0__T_5411_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_5_0__T_5411_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_5_0__T_5411_en = _T_4420 ? 1'h0 : _T_5383;
  assign tensorFile_5_1_rdata_5_addr = tensorFile_5_1_rdata_5_addr_pipe_0;
  assign tensorFile_5_1_rdata_5_data = tensorFile_5_1[tensorFile_5_1_rdata_5_addr]; // @[TensorLoad.scala 222:16:@3455.4]
  assign tensorFile_5_1__T_5411_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_5_1__T_5411_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_5_1__T_5411_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_5_1__T_5411_en = _T_4420 ? 1'h0 : _T_5383;
  assign tensorFile_6_0_rdata_6_addr = tensorFile_6_0_rdata_6_addr_pipe_0;
  assign tensorFile_6_0_rdata_6_data = tensorFile_6_0[tensorFile_6_0_rdata_6_addr]; // @[TensorLoad.scala 222:16:@3456.4]
  assign tensorFile_6_0__T_5498_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_6_0__T_5498_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_6_0__T_5498_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_6_0__T_5498_en = _T_4420 ? 1'h0 : _T_5470;
  assign tensorFile_6_1_rdata_6_addr = tensorFile_6_1_rdata_6_addr_pipe_0;
  assign tensorFile_6_1_rdata_6_data = tensorFile_6_1[tensorFile_6_1_rdata_6_addr]; // @[TensorLoad.scala 222:16:@3456.4]
  assign tensorFile_6_1__T_5498_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_6_1__T_5498_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_6_1__T_5498_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_6_1__T_5498_en = _T_4420 ? 1'h0 : _T_5470;
  assign tensorFile_7_0_rdata_7_addr = tensorFile_7_0_rdata_7_addr_pipe_0;
  assign tensorFile_7_0_rdata_7_data = tensorFile_7_0[tensorFile_7_0_rdata_7_addr]; // @[TensorLoad.scala 222:16:@3457.4]
  assign tensorFile_7_0__T_5585_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_7_0__T_5585_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_7_0__T_5585_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_7_0__T_5585_en = _T_4420 ? 1'h0 : _T_5557;
  assign tensorFile_7_1_rdata_7_addr = tensorFile_7_1_rdata_7_addr_pipe_0;
  assign tensorFile_7_1_rdata_7_data = tensorFile_7_1[tensorFile_7_1_rdata_7_addr]; // @[TensorLoad.scala 222:16:@3457.4]
  assign tensorFile_7_1__T_5585_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_7_1__T_5585_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_7_1__T_5585_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_7_1__T_5585_en = _T_4420 ? 1'h0 : _T_5557;
  assign tensorFile_8_0_rdata_8_addr = tensorFile_8_0_rdata_8_addr_pipe_0;
  assign tensorFile_8_0_rdata_8_data = tensorFile_8_0[tensorFile_8_0_rdata_8_addr]; // @[TensorLoad.scala 222:16:@3458.4]
  assign tensorFile_8_0__T_5672_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_8_0__T_5672_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_8_0__T_5672_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_8_0__T_5672_en = _T_4420 ? 1'h0 : _T_5644;
  assign tensorFile_8_1_rdata_8_addr = tensorFile_8_1_rdata_8_addr_pipe_0;
  assign tensorFile_8_1_rdata_8_data = tensorFile_8_1[tensorFile_8_1_rdata_8_addr]; // @[TensorLoad.scala 222:16:@3458.4]
  assign tensorFile_8_1__T_5672_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_8_1__T_5672_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_8_1__T_5672_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_8_1__T_5672_en = _T_4420 ? 1'h0 : _T_5644;
  assign tensorFile_9_0_rdata_9_addr = tensorFile_9_0_rdata_9_addr_pipe_0;
  assign tensorFile_9_0_rdata_9_data = tensorFile_9_0[tensorFile_9_0_rdata_9_addr]; // @[TensorLoad.scala 222:16:@3459.4]
  assign tensorFile_9_0__T_5759_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_9_0__T_5759_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_9_0__T_5759_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_9_0__T_5759_en = _T_4420 ? 1'h0 : _T_5731;
  assign tensorFile_9_1_rdata_9_addr = tensorFile_9_1_rdata_9_addr_pipe_0;
  assign tensorFile_9_1_rdata_9_data = tensorFile_9_1[tensorFile_9_1_rdata_9_addr]; // @[TensorLoad.scala 222:16:@3459.4]
  assign tensorFile_9_1__T_5759_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_9_1__T_5759_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_9_1__T_5759_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_9_1__T_5759_en = _T_4420 ? 1'h0 : _T_5731;
  assign tensorFile_10_0_rdata_10_addr = tensorFile_10_0_rdata_10_addr_pipe_0;
  assign tensorFile_10_0_rdata_10_data = tensorFile_10_0[tensorFile_10_0_rdata_10_addr]; // @[TensorLoad.scala 222:16:@3460.4]
  assign tensorFile_10_0__T_5846_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_10_0__T_5846_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_10_0__T_5846_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_10_0__T_5846_en = _T_4420 ? 1'h0 : _T_5818;
  assign tensorFile_10_1_rdata_10_addr = tensorFile_10_1_rdata_10_addr_pipe_0;
  assign tensorFile_10_1_rdata_10_data = tensorFile_10_1[tensorFile_10_1_rdata_10_addr]; // @[TensorLoad.scala 222:16:@3460.4]
  assign tensorFile_10_1__T_5846_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_10_1__T_5846_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_10_1__T_5846_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_10_1__T_5846_en = _T_4420 ? 1'h0 : _T_5818;
  assign tensorFile_11_0_rdata_11_addr = tensorFile_11_0_rdata_11_addr_pipe_0;
  assign tensorFile_11_0_rdata_11_data = tensorFile_11_0[tensorFile_11_0_rdata_11_addr]; // @[TensorLoad.scala 222:16:@3461.4]
  assign tensorFile_11_0__T_5933_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_11_0__T_5933_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_11_0__T_5933_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_11_0__T_5933_en = _T_4420 ? 1'h0 : _T_5905;
  assign tensorFile_11_1_rdata_11_addr = tensorFile_11_1_rdata_11_addr_pipe_0;
  assign tensorFile_11_1_rdata_11_data = tensorFile_11_1[tensorFile_11_1_rdata_11_addr]; // @[TensorLoad.scala 222:16:@3461.4]
  assign tensorFile_11_1__T_5933_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_11_1__T_5933_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_11_1__T_5933_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_11_1__T_5933_en = _T_4420 ? 1'h0 : _T_5905;
  assign tensorFile_12_0_rdata_12_addr = tensorFile_12_0_rdata_12_addr_pipe_0;
  assign tensorFile_12_0_rdata_12_data = tensorFile_12_0[tensorFile_12_0_rdata_12_addr]; // @[TensorLoad.scala 222:16:@3462.4]
  assign tensorFile_12_0__T_6020_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_12_0__T_6020_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_12_0__T_6020_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_12_0__T_6020_en = _T_4420 ? 1'h0 : _T_5992;
  assign tensorFile_12_1_rdata_12_addr = tensorFile_12_1_rdata_12_addr_pipe_0;
  assign tensorFile_12_1_rdata_12_data = tensorFile_12_1[tensorFile_12_1_rdata_12_addr]; // @[TensorLoad.scala 222:16:@3462.4]
  assign tensorFile_12_1__T_6020_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_12_1__T_6020_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_12_1__T_6020_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_12_1__T_6020_en = _T_4420 ? 1'h0 : _T_5992;
  assign tensorFile_13_0_rdata_13_addr = tensorFile_13_0_rdata_13_addr_pipe_0;
  assign tensorFile_13_0_rdata_13_data = tensorFile_13_0[tensorFile_13_0_rdata_13_addr]; // @[TensorLoad.scala 222:16:@3463.4]
  assign tensorFile_13_0__T_6107_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_13_0__T_6107_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_13_0__T_6107_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_13_0__T_6107_en = _T_4420 ? 1'h0 : _T_6079;
  assign tensorFile_13_1_rdata_13_addr = tensorFile_13_1_rdata_13_addr_pipe_0;
  assign tensorFile_13_1_rdata_13_data = tensorFile_13_1[tensorFile_13_1_rdata_13_addr]; // @[TensorLoad.scala 222:16:@3463.4]
  assign tensorFile_13_1__T_6107_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_13_1__T_6107_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_13_1__T_6107_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_13_1__T_6107_en = _T_4420 ? 1'h0 : _T_6079;
  assign tensorFile_14_0_rdata_14_addr = tensorFile_14_0_rdata_14_addr_pipe_0;
  assign tensorFile_14_0_rdata_14_data = tensorFile_14_0[tensorFile_14_0_rdata_14_addr]; // @[TensorLoad.scala 222:16:@3464.4]
  assign tensorFile_14_0__T_6194_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_14_0__T_6194_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_14_0__T_6194_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_14_0__T_6194_en = _T_4420 ? 1'h0 : _T_6166;
  assign tensorFile_14_1_rdata_14_addr = tensorFile_14_1_rdata_14_addr_pipe_0;
  assign tensorFile_14_1_rdata_14_data = tensorFile_14_1[tensorFile_14_1_rdata_14_addr]; // @[TensorLoad.scala 222:16:@3464.4]
  assign tensorFile_14_1__T_6194_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_14_1__T_6194_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_14_1__T_6194_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_14_1__T_6194_en = _T_4420 ? 1'h0 : _T_6166;
  assign tensorFile_15_0_rdata_15_addr = tensorFile_15_0_rdata_15_addr_pipe_0;
  assign tensorFile_15_0_rdata_15_data = tensorFile_15_0[tensorFile_15_0_rdata_15_addr]; // @[TensorLoad.scala 222:16:@3465.4]
  assign tensorFile_15_0__T_6281_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_15_0__T_6281_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_15_0__T_6281_mask = _T_4420 ? 1'h1 : wmask_0_0;
  assign tensorFile_15_0__T_6281_en = _T_4420 ? 1'h0 : _T_4523;
  assign tensorFile_15_1_rdata_15_addr = tensorFile_15_1_rdata_15_addr_pipe_0;
  assign tensorFile_15_1_rdata_15_data = tensorFile_15_1[tensorFile_15_1_rdata_15_addr]; // @[TensorLoad.scala 222:16:@3465.4]
  assign tensorFile_15_1__T_6281_data = _T_4420 ? 64'h0 : wdata_0_0;
  assign tensorFile_15_1__T_6281_addr = _T_4420 ? 10'h0 : waddr_cur;
  assign tensorFile_15_1__T_6281_mask = _T_4420 ? 1'h1 : tag;
  assign tensorFile_15_1__T_6281_en = _T_4420 ? 1'h0 : _T_4523;
  assign dec_sram_offset = io_inst[24:9]; // @[TensorLoad.scala 51:29:@3147.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorLoad.scala 51:29:@3155.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorLoad.scala 51:29:@3159.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorLoad.scala 51:29:@3161.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorLoad.scala 51:29:@3163.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorLoad.scala 51:29:@3165.4]
  assign _T_4394 = 3'h0 == state; // @[Conditional.scala 37:30:@3186.4]
  assign _T_4396 = dec_ypad_0 != 4'h0; // @[TensorLoad.scala 71:25:@3189.8]
  assign _T_4398 = dec_xpad_0 != 4'h0; // @[TensorLoad.scala 73:31:@3194.10]
  assign _GEN_0 = _T_4398 ? 3'h2 : 3'h3; // @[TensorLoad.scala 73:40:@3195.10]
  assign _GEN_1 = _T_4396 ? 3'h1 : _GEN_0; // @[TensorLoad.scala 71:34:@3190.8]
  assign _GEN_2 = io_start ? _GEN_1 : state; // @[TensorLoad.scala 70:22:@3188.6]
  assign _T_4399 = 3'h1 == state; // @[Conditional.scala 37:30:@3204.6]
  assign _GEN_4 = yPadCtrl0_io_done ? _GEN_0 : state; // @[TensorLoad.scala 81:31:@3206.8]
  assign _T_4402 = 3'h2 == state; // @[Conditional.scala 37:30:@3217.8]
  assign _GEN_5 = xPadCtrl0_io_done ? 3'h3 : state; // @[TensorLoad.scala 90:31:@3219.10]
  assign _T_4403 = 3'h3 == state; // @[Conditional.scala 37:30:@3224.10]
  assign _GEN_6 = io_vme_rd_cmd_ready ? 3'h4 : state; // @[TensorLoad.scala 95:33:@3226.12]
  assign _T_4404 = 3'h4 == state; // @[Conditional.scala 37:30:@3231.12]
  assign _T_4406 = dec_xpad_1 != 4'h0; // @[TensorLoad.scala 102:27:@3235.18]
  assign _T_4408 = dec_ypad_1 != 4'h0; // @[TensorLoad.scala 104:33:@3240.20]
  assign _GEN_7 = _T_4408 ? 3'h6 : 3'h0; // @[TensorLoad.scala 104:42:@3241.20]
  assign _GEN_8 = _T_4406 ? 3'h5 : _GEN_7; // @[TensorLoad.scala 102:36:@3236.18]
  assign _GEN_10 = _T_4406 ? 3'h5 : _GEN_0; // @[TensorLoad.scala 110:36:@3251.20]
  assign _GEN_11 = dataCtrl_io_split ? 3'h3 : state; // @[TensorLoad.scala 117:39:@3264.20]
  assign _GEN_12 = dataCtrl_io_stride ? _GEN_10 : _GEN_11; // @[TensorLoad.scala 109:40:@3249.18]
  assign _GEN_13 = dataCtrl_io_done ? _GEN_8 : _GEN_12; // @[TensorLoad.scala 101:32:@3234.16]
  assign _GEN_14 = io_vme_rd_data_valid ? _GEN_13 : state; // @[TensorLoad.scala 100:34:@3233.14]
  assign _T_4413 = 3'h5 == state; // @[Conditional.scala 37:30:@3270.14]
  assign _GEN_17 = dataCtrlDone ? _GEN_7 : _GEN_0; // @[TensorLoad.scala 124:28:@3273.18]
  assign _GEN_18 = xPadCtrl1_io_done ? _GEN_17 : state; // @[TensorLoad.scala 123:31:@3272.16]
  assign _T_4418 = 3'h6 == state; // @[Conditional.scala 37:30:@3294.16]
  assign _T_4419 = yPadCtrl1_io_done & dataCtrlDone; // @[TensorLoad.scala 140:30:@3296.18]
  assign _GEN_19 = _T_4419 ? 3'h0 : state; // @[TensorLoad.scala 140:47:@3297.18]
  assign _GEN_20 = _T_4418 ? _GEN_19 : state; // @[Conditional.scala 39:67:@3295.16]
  assign _GEN_21 = _T_4413 ? _GEN_18 : _GEN_20; // @[Conditional.scala 39:67:@3271.14]
  assign _GEN_22 = _T_4404 ? _GEN_14 : _GEN_21; // @[Conditional.scala 39:67:@3232.12]
  assign _GEN_23 = _T_4403 ? _GEN_6 : _GEN_22; // @[Conditional.scala 39:67:@3225.10]
  assign _GEN_24 = _T_4402 ? _GEN_5 : _GEN_23; // @[Conditional.scala 39:67:@3218.8]
  assign _GEN_25 = _T_4399 ? _GEN_4 : _GEN_24; // @[Conditional.scala 39:67:@3205.6]
  assign _GEN_26 = _T_4394 ? _GEN_2 : _GEN_25; // @[Conditional.scala 40:58:@3187.4]
  assign _T_4420 = state == 3'h0; // @[TensorLoad.scala 147:30:@3301.4]
  assign _T_4421 = _T_4420 & io_start; // @[TensorLoad.scala 147:40:@3302.4]
  assign _T_4423 = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[Decoupled.scala 37:37:@3308.4]
  assign _T_4428 = _T_4423 & dataCtrl_io_done; // @[TensorLoad.scala 156:36:@3318.6]
  assign _GEN_27 = _T_4428 ? 1'h1 : dataCtrlDone; // @[TensorLoad.scala 156:57:@3319.6]
  assign _GEN_28 = _T_4420 ? 1'h0 : _GEN_27; // @[TensorLoad.scala 154:25:@3313.4]
  assign _T_4433 = _T_4396 & _T_4420; // @[TensorLoad.scala 161:44:@3324.4]
  assign _T_4440 = dec_xpad_1 == 4'h0; // @[TensorLoad.scala 164:61:@3330.4]
  assign _T_4441 = _T_4428 & _T_4440; // @[TensorLoad.scala 164:48:@3331.4]
  assign _T_4442 = state == 3'h5; // @[TensorLoad.scala 165:14:@3332.4]
  assign _T_4443 = _T_4442 & xPadCtrl1_io_done; // @[TensorLoad.scala 165:25:@3333.4]
  assign _T_4444 = _T_4443 & dataCtrlDone; // @[TensorLoad.scala 165:45:@3334.4]
  assign _T_4445 = _T_4441 | _T_4444; // @[TensorLoad.scala 164:70:@3335.4]
  assign _T_4451 = state == 3'h1; // @[TensorLoad.scala 169:14:@3341.4]
  assign _T_4452 = _T_4451 & yPadCtrl0_io_done; // @[TensorLoad.scala 169:25:@3342.4]
  assign _T_4453 = _T_4421 | _T_4452; // @[TensorLoad.scala 168:35:@3343.4]
  assign _T_4455 = ~ dataCtrlDone; // @[TensorLoad.scala 170:32:@3345.4]
  assign _T_4456 = _T_4423 & _T_4455; // @[TensorLoad.scala 170:30:@3346.4]
  assign _T_4457 = _T_4456 & dataCtrl_io_stride; // @[TensorLoad.scala 170:46:@3347.4]
  assign _T_4460 = _T_4457 & _T_4440; // @[TensorLoad.scala 170:67:@3349.4]
  assign _T_4461 = _T_4453 | _T_4460; // @[TensorLoad.scala 169:46:@3350.4]
  assign _T_4465 = _T_4443 & _T_4455; // @[TensorLoad.scala 171:45:@3354.4]
  assign _T_4466 = _T_4461 | _T_4465; // @[TensorLoad.scala 170:89:@3355.4]
  assign _T_4471 = _T_4406 & _T_4423; // @[TensorLoad.scala 173:44:@3360.4]
  assign _T_4472 = ~ dataCtrl_io_done; // @[TensorLoad.scala 174:28:@3361.4]
  assign _T_4473 = _T_4472 & dataCtrl_io_stride; // @[TensorLoad.scala 174:46:@3362.4]
  assign _T_4476 = _T_4473 & _T_4406; // @[TensorLoad.scala 174:67:@3364.4]
  assign _T_4477 = dataCtrl_io_done | _T_4476; // @[TensorLoad.scala 174:25:@3365.4]
  assign _T_4479 = state == 3'h3; // @[TensorLoad.scala 182:32:@3372.4]
  assign _T_4482 = state == 3'h2; // @[TensorLoad.scala 190:11:@3379.4]
  assign _T_4483 = _T_4451 | _T_4482; // @[TensorLoad.scala 189:36:@3380.4]
  assign _T_4485 = _T_4483 | _T_4442; // @[TensorLoad.scala 190:22:@3382.4]
  assign _T_4486 = state == 3'h6; // @[TensorLoad.scala 192:11:@3383.4]
  assign isZeroPad = _T_4485 | _T_4486; // @[TensorLoad.scala 191:22:@3384.4]
  assign _T_4489 = _T_4420 | _T_4479; // @[TensorLoad.scala 194:24:@3387.4]
  assign _T_4492 = _T_4489 | tag; // @[TensorLoad.scala 194:46:@3389.4]
  assign _T_4495 = _T_4423 | isZeroPad; // @[TensorLoad.scala 196:36:@3395.6]
  assign _T_4497 = tag + 1'h1; // @[TensorLoad.scala 197:16:@3397.8]
  assign _T_4498 = tag + 1'h1; // @[TensorLoad.scala 197:16:@3398.8]
  assign _GEN_29 = _T_4495 ? _T_4498 : tag; // @[TensorLoad.scala 196:50:@3396.6]
  assign _T_4500 = _T_4420 | dataCtrlDone; // @[TensorLoad.scala 200:24:@3402.4]
  assign _T_4502 = set == 4'hf; // @[TensorLoad.scala 200:48:@3403.4]
  assign _T_4505 = _T_4502 & tag; // @[TensorLoad.scala 200:76:@3405.4]
  assign _T_4506 = _T_4500 | _T_4505; // @[TensorLoad.scala 200:40:@3406.4]
  assign _T_4512 = _T_4495 & tag; // @[TensorLoad.scala 202:51:@3414.6]
  assign _T_4514 = set + 4'h1; // @[TensorLoad.scala 203:16:@3416.8]
  assign _T_4515 = set + 4'h1; // @[TensorLoad.scala 203:16:@3417.8]
  assign _GEN_31 = _T_4512 ? _T_4515 : set; // @[TensorLoad.scala 202:86:@3415.6]
  assign _T_4523 = _T_4495 & _T_4502; // @[TensorLoad.scala 212:5:@3431.6]
  assign _T_4526 = _T_4523 & tag; // @[TensorLoad.scala 213:5:@3433.6]
  assign _T_4528 = waddr_cur + 10'h1; // @[TensorLoad.scala 215:28:@3435.8]
  assign _T_4529 = waddr_cur + 10'h1; // @[TensorLoad.scala 215:28:@3436.8]
  assign _T_4531 = dataCtrl_io_stride & _T_4423; // @[TensorLoad.scala 216:33:@3441.8]
  assign _GEN_426 = {{6'd0}, waddr_nxt}; // @[TensorLoad.scala 217:28:@3443.10]
  assign _T_4532 = _GEN_426 + dec_xsize; // @[TensorLoad.scala 217:28:@3443.10]
  assign _T_4533 = _GEN_426 + dec_xsize; // @[TensorLoad.scala 217:28:@3444.10]
  assign _GEN_33 = _T_4531 ? _T_4533 : {{6'd0}, waddr_cur}; // @[TensorLoad.scala 216:59:@3442.8]
  assign _GEN_34 = _T_4531 ? _T_4533 : {{6'd0}, waddr_nxt}; // @[TensorLoad.scala 216:59:@3442.8]
  assign _GEN_35 = _T_4526 ? {{6'd0}, _T_4529} : _GEN_33; // @[TensorLoad.scala 214:3:@3434.6]
  assign _GEN_36 = _T_4526 ? {{6'd0}, waddr_nxt} : _GEN_34; // @[TensorLoad.scala 214:3:@3434.6]
  assign _GEN_37 = _T_4420 ? dec_sram_offset : _GEN_35; // @[TensorLoad.scala 208:25:@3423.4]
  assign _GEN_38 = _T_4420 ? dec_sram_offset : _GEN_36; // @[TensorLoad.scala 208:25:@3423.4]
  assign wmask_0_0 = tag == 1'h0; // @[TensorLoad.scala 235:26:@3501.4]
  assign wdata_0_0 = isZeroPad ? 64'h0 : io_vme_rd_data_bits; // @[TensorLoad.scala 236:25:@3503.4]
  assign _T_4947 = set == 4'h0; // @[TensorLoad.scala 242:51:@3534.4]
  assign _T_4948 = _T_4495 & _T_4947; // @[TensorLoad.scala 242:45:@3535.4]
  assign _T_5034 = set == 4'h1; // @[TensorLoad.scala 242:51:@3585.4]
  assign _T_5035 = _T_4495 & _T_5034; // @[TensorLoad.scala 242:45:@3586.4]
  assign _T_5121 = set == 4'h2; // @[TensorLoad.scala 242:51:@3636.4]
  assign _T_5122 = _T_4495 & _T_5121; // @[TensorLoad.scala 242:45:@3637.4]
  assign _T_5208 = set == 4'h3; // @[TensorLoad.scala 242:51:@3687.4]
  assign _T_5209 = _T_4495 & _T_5208; // @[TensorLoad.scala 242:45:@3688.4]
  assign _T_5295 = set == 4'h4; // @[TensorLoad.scala 242:51:@3738.4]
  assign _T_5296 = _T_4495 & _T_5295; // @[TensorLoad.scala 242:45:@3739.4]
  assign _T_5382 = set == 4'h5; // @[TensorLoad.scala 242:51:@3789.4]
  assign _T_5383 = _T_4495 & _T_5382; // @[TensorLoad.scala 242:45:@3790.4]
  assign _T_5469 = set == 4'h6; // @[TensorLoad.scala 242:51:@3840.4]
  assign _T_5470 = _T_4495 & _T_5469; // @[TensorLoad.scala 242:45:@3841.4]
  assign _T_5556 = set == 4'h7; // @[TensorLoad.scala 242:51:@3891.4]
  assign _T_5557 = _T_4495 & _T_5556; // @[TensorLoad.scala 242:45:@3892.4]
  assign _T_5643 = set == 4'h8; // @[TensorLoad.scala 242:51:@3942.4]
  assign _T_5644 = _T_4495 & _T_5643; // @[TensorLoad.scala 242:45:@3943.4]
  assign _T_5730 = set == 4'h9; // @[TensorLoad.scala 242:51:@3993.4]
  assign _T_5731 = _T_4495 & _T_5730; // @[TensorLoad.scala 242:45:@3994.4]
  assign _T_5817 = set == 4'ha; // @[TensorLoad.scala 242:51:@4044.4]
  assign _T_5818 = _T_4495 & _T_5817; // @[TensorLoad.scala 242:45:@4045.4]
  assign _T_5904 = set == 4'hb; // @[TensorLoad.scala 242:51:@4095.4]
  assign _T_5905 = _T_4495 & _T_5904; // @[TensorLoad.scala 242:45:@4096.4]
  assign _T_5991 = set == 4'hc; // @[TensorLoad.scala 242:51:@4146.4]
  assign _T_5992 = _T_4495 & _T_5991; // @[TensorLoad.scala 242:45:@4147.4]
  assign _T_6078 = set == 4'hd; // @[TensorLoad.scala 242:51:@4197.4]
  assign _T_6079 = _T_4495 & _T_6078; // @[TensorLoad.scala 242:45:@4198.4]
  assign _T_6165 = set == 4'he; // @[TensorLoad.scala 242:51:@4248.4]
  assign _T_6166 = _T_4495 & _T_6165; // @[TensorLoad.scala 242:45:@4249.4]
  assign _GEN_216 = io_tensor_rd_idx_valid; // @[TensorLoad.scala 256:26:@4322.4]
  assign _T_6482 = {tensorFile_0_1_rdata_0_data,tensorFile_0_0_rdata_0_data}; // @[TensorLoad.scala 259:38:@4448.4]
  assign _T_6624 = {tensorFile_1_1_rdata_1_data,tensorFile_1_0_rdata_1_data}; // @[TensorLoad.scala 259:38:@4500.4]
  assign _T_6766 = {tensorFile_2_1_rdata_2_data,tensorFile_2_0_rdata_2_data}; // @[TensorLoad.scala 259:38:@4552.4]
  assign _T_6908 = {tensorFile_3_1_rdata_3_data,tensorFile_3_0_rdata_3_data}; // @[TensorLoad.scala 259:38:@4604.4]
  assign _T_7050 = {tensorFile_4_1_rdata_4_data,tensorFile_4_0_rdata_4_data}; // @[TensorLoad.scala 259:38:@4656.4]
  assign _T_7192 = {tensorFile_5_1_rdata_5_data,tensorFile_5_0_rdata_5_data}; // @[TensorLoad.scala 259:38:@4708.4]
  assign _T_7334 = {tensorFile_6_1_rdata_6_data,tensorFile_6_0_rdata_6_data}; // @[TensorLoad.scala 259:38:@4760.4]
  assign _T_7476 = {tensorFile_7_1_rdata_7_data,tensorFile_7_0_rdata_7_data}; // @[TensorLoad.scala 259:38:@4812.4]
  assign _T_7618 = {tensorFile_8_1_rdata_8_data,tensorFile_8_0_rdata_8_data}; // @[TensorLoad.scala 259:38:@4864.4]
  assign _T_7760 = {tensorFile_9_1_rdata_9_data,tensorFile_9_0_rdata_9_data}; // @[TensorLoad.scala 259:38:@4916.4]
  assign _T_7902 = {tensorFile_10_1_rdata_10_data,tensorFile_10_0_rdata_10_data}; // @[TensorLoad.scala 259:38:@4968.4]
  assign _T_8044 = {tensorFile_11_1_rdata_11_data,tensorFile_11_0_rdata_11_data}; // @[TensorLoad.scala 259:38:@5020.4]
  assign _T_8186 = {tensorFile_12_1_rdata_12_data,tensorFile_12_0_rdata_12_data}; // @[TensorLoad.scala 259:38:@5072.4]
  assign _T_8328 = {tensorFile_13_1_rdata_13_data,tensorFile_13_0_rdata_13_data}; // @[TensorLoad.scala 259:38:@5124.4]
  assign _T_8470 = {tensorFile_14_1_rdata_14_data,tensorFile_14_0_rdata_14_data}; // @[TensorLoad.scala 259:38:@5176.4]
  assign _T_8612 = {tensorFile_15_1_rdata_15_data,tensorFile_15_0_rdata_15_data}; // @[TensorLoad.scala 259:38:@5228.4]
  assign _T_8760 = dec_ypad_1 == 4'h0; // @[TensorLoad.scala 263:96:@5284.4]
  assign done_no_pad = _T_4441 & _T_8760; // @[TensorLoad.scala 263:83:@5285.4]
  assign done_x_pad = _T_4444 & _T_8760; // @[TensorLoad.scala 264:72:@5290.4]
  assign _T_8767 = _T_4486 & dataCtrlDone; // @[TensorLoad.scala 265:37:@5292.4]
  assign done_y_pad = _T_8767 & yPadCtrl1_io_done; // @[TensorLoad.scala 265:52:@5293.4]
  assign _T_8768 = done_no_pad | done_x_pad; // @[TensorLoad.scala 266:26:@5294.4]
  assign io_done = _T_8768 | done_y_pad; // @[TensorLoad.scala 266:11:@5296.4]
  assign io_vme_rd_cmd_valid = state == 3'h3; // @[TensorLoad.scala 182:23:@3373.4]
  assign io_vme_rd_cmd_bits_addr = dataCtrl_io_addr; // @[TensorLoad.scala 183:27:@3374.4]
  assign io_vme_rd_cmd_bits_len = dataCtrl_io_len; // @[TensorLoad.scala 184:26:@3375.4]
  assign io_vme_rd_data_ready = state == 3'h4; // @[TensorLoad.scala 186:24:@3377.4]
  assign io_tensor_rd_data_valid = rvalid; // @[TensorLoad.scala 253:27:@4319.4]
  assign io_tensor_rd_data_bits_0_0 = _T_6482[7:0]; // @[TensorLoad.scala 259:33:@4484.4]
  assign io_tensor_rd_data_bits_0_1 = _T_6482[15:8]; // @[TensorLoad.scala 259:33:@4485.4]
  assign io_tensor_rd_data_bits_0_2 = _T_6482[23:16]; // @[TensorLoad.scala 259:33:@4486.4]
  assign io_tensor_rd_data_bits_0_3 = _T_6482[31:24]; // @[TensorLoad.scala 259:33:@4487.4]
  assign io_tensor_rd_data_bits_0_4 = _T_6482[39:32]; // @[TensorLoad.scala 259:33:@4488.4]
  assign io_tensor_rd_data_bits_0_5 = _T_6482[47:40]; // @[TensorLoad.scala 259:33:@4489.4]
  assign io_tensor_rd_data_bits_0_6 = _T_6482[55:48]; // @[TensorLoad.scala 259:33:@4490.4]
  assign io_tensor_rd_data_bits_0_7 = _T_6482[63:56]; // @[TensorLoad.scala 259:33:@4491.4]
  assign io_tensor_rd_data_bits_0_8 = _T_6482[71:64]; // @[TensorLoad.scala 259:33:@4492.4]
  assign io_tensor_rd_data_bits_0_9 = _T_6482[79:72]; // @[TensorLoad.scala 259:33:@4493.4]
  assign io_tensor_rd_data_bits_0_10 = _T_6482[87:80]; // @[TensorLoad.scala 259:33:@4494.4]
  assign io_tensor_rd_data_bits_0_11 = _T_6482[95:88]; // @[TensorLoad.scala 259:33:@4495.4]
  assign io_tensor_rd_data_bits_0_12 = _T_6482[103:96]; // @[TensorLoad.scala 259:33:@4496.4]
  assign io_tensor_rd_data_bits_0_13 = _T_6482[111:104]; // @[TensorLoad.scala 259:33:@4497.4]
  assign io_tensor_rd_data_bits_0_14 = _T_6482[119:112]; // @[TensorLoad.scala 259:33:@4498.4]
  assign io_tensor_rd_data_bits_0_15 = _T_6482[127:120]; // @[TensorLoad.scala 259:33:@4499.4]
  assign io_tensor_rd_data_bits_1_0 = _T_6624[7:0]; // @[TensorLoad.scala 259:33:@4536.4]
  assign io_tensor_rd_data_bits_1_1 = _T_6624[15:8]; // @[TensorLoad.scala 259:33:@4537.4]
  assign io_tensor_rd_data_bits_1_2 = _T_6624[23:16]; // @[TensorLoad.scala 259:33:@4538.4]
  assign io_tensor_rd_data_bits_1_3 = _T_6624[31:24]; // @[TensorLoad.scala 259:33:@4539.4]
  assign io_tensor_rd_data_bits_1_4 = _T_6624[39:32]; // @[TensorLoad.scala 259:33:@4540.4]
  assign io_tensor_rd_data_bits_1_5 = _T_6624[47:40]; // @[TensorLoad.scala 259:33:@4541.4]
  assign io_tensor_rd_data_bits_1_6 = _T_6624[55:48]; // @[TensorLoad.scala 259:33:@4542.4]
  assign io_tensor_rd_data_bits_1_7 = _T_6624[63:56]; // @[TensorLoad.scala 259:33:@4543.4]
  assign io_tensor_rd_data_bits_1_8 = _T_6624[71:64]; // @[TensorLoad.scala 259:33:@4544.4]
  assign io_tensor_rd_data_bits_1_9 = _T_6624[79:72]; // @[TensorLoad.scala 259:33:@4545.4]
  assign io_tensor_rd_data_bits_1_10 = _T_6624[87:80]; // @[TensorLoad.scala 259:33:@4546.4]
  assign io_tensor_rd_data_bits_1_11 = _T_6624[95:88]; // @[TensorLoad.scala 259:33:@4547.4]
  assign io_tensor_rd_data_bits_1_12 = _T_6624[103:96]; // @[TensorLoad.scala 259:33:@4548.4]
  assign io_tensor_rd_data_bits_1_13 = _T_6624[111:104]; // @[TensorLoad.scala 259:33:@4549.4]
  assign io_tensor_rd_data_bits_1_14 = _T_6624[119:112]; // @[TensorLoad.scala 259:33:@4550.4]
  assign io_tensor_rd_data_bits_1_15 = _T_6624[127:120]; // @[TensorLoad.scala 259:33:@4551.4]
  assign io_tensor_rd_data_bits_2_0 = _T_6766[7:0]; // @[TensorLoad.scala 259:33:@4588.4]
  assign io_tensor_rd_data_bits_2_1 = _T_6766[15:8]; // @[TensorLoad.scala 259:33:@4589.4]
  assign io_tensor_rd_data_bits_2_2 = _T_6766[23:16]; // @[TensorLoad.scala 259:33:@4590.4]
  assign io_tensor_rd_data_bits_2_3 = _T_6766[31:24]; // @[TensorLoad.scala 259:33:@4591.4]
  assign io_tensor_rd_data_bits_2_4 = _T_6766[39:32]; // @[TensorLoad.scala 259:33:@4592.4]
  assign io_tensor_rd_data_bits_2_5 = _T_6766[47:40]; // @[TensorLoad.scala 259:33:@4593.4]
  assign io_tensor_rd_data_bits_2_6 = _T_6766[55:48]; // @[TensorLoad.scala 259:33:@4594.4]
  assign io_tensor_rd_data_bits_2_7 = _T_6766[63:56]; // @[TensorLoad.scala 259:33:@4595.4]
  assign io_tensor_rd_data_bits_2_8 = _T_6766[71:64]; // @[TensorLoad.scala 259:33:@4596.4]
  assign io_tensor_rd_data_bits_2_9 = _T_6766[79:72]; // @[TensorLoad.scala 259:33:@4597.4]
  assign io_tensor_rd_data_bits_2_10 = _T_6766[87:80]; // @[TensorLoad.scala 259:33:@4598.4]
  assign io_tensor_rd_data_bits_2_11 = _T_6766[95:88]; // @[TensorLoad.scala 259:33:@4599.4]
  assign io_tensor_rd_data_bits_2_12 = _T_6766[103:96]; // @[TensorLoad.scala 259:33:@4600.4]
  assign io_tensor_rd_data_bits_2_13 = _T_6766[111:104]; // @[TensorLoad.scala 259:33:@4601.4]
  assign io_tensor_rd_data_bits_2_14 = _T_6766[119:112]; // @[TensorLoad.scala 259:33:@4602.4]
  assign io_tensor_rd_data_bits_2_15 = _T_6766[127:120]; // @[TensorLoad.scala 259:33:@4603.4]
  assign io_tensor_rd_data_bits_3_0 = _T_6908[7:0]; // @[TensorLoad.scala 259:33:@4640.4]
  assign io_tensor_rd_data_bits_3_1 = _T_6908[15:8]; // @[TensorLoad.scala 259:33:@4641.4]
  assign io_tensor_rd_data_bits_3_2 = _T_6908[23:16]; // @[TensorLoad.scala 259:33:@4642.4]
  assign io_tensor_rd_data_bits_3_3 = _T_6908[31:24]; // @[TensorLoad.scala 259:33:@4643.4]
  assign io_tensor_rd_data_bits_3_4 = _T_6908[39:32]; // @[TensorLoad.scala 259:33:@4644.4]
  assign io_tensor_rd_data_bits_3_5 = _T_6908[47:40]; // @[TensorLoad.scala 259:33:@4645.4]
  assign io_tensor_rd_data_bits_3_6 = _T_6908[55:48]; // @[TensorLoad.scala 259:33:@4646.4]
  assign io_tensor_rd_data_bits_3_7 = _T_6908[63:56]; // @[TensorLoad.scala 259:33:@4647.4]
  assign io_tensor_rd_data_bits_3_8 = _T_6908[71:64]; // @[TensorLoad.scala 259:33:@4648.4]
  assign io_tensor_rd_data_bits_3_9 = _T_6908[79:72]; // @[TensorLoad.scala 259:33:@4649.4]
  assign io_tensor_rd_data_bits_3_10 = _T_6908[87:80]; // @[TensorLoad.scala 259:33:@4650.4]
  assign io_tensor_rd_data_bits_3_11 = _T_6908[95:88]; // @[TensorLoad.scala 259:33:@4651.4]
  assign io_tensor_rd_data_bits_3_12 = _T_6908[103:96]; // @[TensorLoad.scala 259:33:@4652.4]
  assign io_tensor_rd_data_bits_3_13 = _T_6908[111:104]; // @[TensorLoad.scala 259:33:@4653.4]
  assign io_tensor_rd_data_bits_3_14 = _T_6908[119:112]; // @[TensorLoad.scala 259:33:@4654.4]
  assign io_tensor_rd_data_bits_3_15 = _T_6908[127:120]; // @[TensorLoad.scala 259:33:@4655.4]
  assign io_tensor_rd_data_bits_4_0 = _T_7050[7:0]; // @[TensorLoad.scala 259:33:@4692.4]
  assign io_tensor_rd_data_bits_4_1 = _T_7050[15:8]; // @[TensorLoad.scala 259:33:@4693.4]
  assign io_tensor_rd_data_bits_4_2 = _T_7050[23:16]; // @[TensorLoad.scala 259:33:@4694.4]
  assign io_tensor_rd_data_bits_4_3 = _T_7050[31:24]; // @[TensorLoad.scala 259:33:@4695.4]
  assign io_tensor_rd_data_bits_4_4 = _T_7050[39:32]; // @[TensorLoad.scala 259:33:@4696.4]
  assign io_tensor_rd_data_bits_4_5 = _T_7050[47:40]; // @[TensorLoad.scala 259:33:@4697.4]
  assign io_tensor_rd_data_bits_4_6 = _T_7050[55:48]; // @[TensorLoad.scala 259:33:@4698.4]
  assign io_tensor_rd_data_bits_4_7 = _T_7050[63:56]; // @[TensorLoad.scala 259:33:@4699.4]
  assign io_tensor_rd_data_bits_4_8 = _T_7050[71:64]; // @[TensorLoad.scala 259:33:@4700.4]
  assign io_tensor_rd_data_bits_4_9 = _T_7050[79:72]; // @[TensorLoad.scala 259:33:@4701.4]
  assign io_tensor_rd_data_bits_4_10 = _T_7050[87:80]; // @[TensorLoad.scala 259:33:@4702.4]
  assign io_tensor_rd_data_bits_4_11 = _T_7050[95:88]; // @[TensorLoad.scala 259:33:@4703.4]
  assign io_tensor_rd_data_bits_4_12 = _T_7050[103:96]; // @[TensorLoad.scala 259:33:@4704.4]
  assign io_tensor_rd_data_bits_4_13 = _T_7050[111:104]; // @[TensorLoad.scala 259:33:@4705.4]
  assign io_tensor_rd_data_bits_4_14 = _T_7050[119:112]; // @[TensorLoad.scala 259:33:@4706.4]
  assign io_tensor_rd_data_bits_4_15 = _T_7050[127:120]; // @[TensorLoad.scala 259:33:@4707.4]
  assign io_tensor_rd_data_bits_5_0 = _T_7192[7:0]; // @[TensorLoad.scala 259:33:@4744.4]
  assign io_tensor_rd_data_bits_5_1 = _T_7192[15:8]; // @[TensorLoad.scala 259:33:@4745.4]
  assign io_tensor_rd_data_bits_5_2 = _T_7192[23:16]; // @[TensorLoad.scala 259:33:@4746.4]
  assign io_tensor_rd_data_bits_5_3 = _T_7192[31:24]; // @[TensorLoad.scala 259:33:@4747.4]
  assign io_tensor_rd_data_bits_5_4 = _T_7192[39:32]; // @[TensorLoad.scala 259:33:@4748.4]
  assign io_tensor_rd_data_bits_5_5 = _T_7192[47:40]; // @[TensorLoad.scala 259:33:@4749.4]
  assign io_tensor_rd_data_bits_5_6 = _T_7192[55:48]; // @[TensorLoad.scala 259:33:@4750.4]
  assign io_tensor_rd_data_bits_5_7 = _T_7192[63:56]; // @[TensorLoad.scala 259:33:@4751.4]
  assign io_tensor_rd_data_bits_5_8 = _T_7192[71:64]; // @[TensorLoad.scala 259:33:@4752.4]
  assign io_tensor_rd_data_bits_5_9 = _T_7192[79:72]; // @[TensorLoad.scala 259:33:@4753.4]
  assign io_tensor_rd_data_bits_5_10 = _T_7192[87:80]; // @[TensorLoad.scala 259:33:@4754.4]
  assign io_tensor_rd_data_bits_5_11 = _T_7192[95:88]; // @[TensorLoad.scala 259:33:@4755.4]
  assign io_tensor_rd_data_bits_5_12 = _T_7192[103:96]; // @[TensorLoad.scala 259:33:@4756.4]
  assign io_tensor_rd_data_bits_5_13 = _T_7192[111:104]; // @[TensorLoad.scala 259:33:@4757.4]
  assign io_tensor_rd_data_bits_5_14 = _T_7192[119:112]; // @[TensorLoad.scala 259:33:@4758.4]
  assign io_tensor_rd_data_bits_5_15 = _T_7192[127:120]; // @[TensorLoad.scala 259:33:@4759.4]
  assign io_tensor_rd_data_bits_6_0 = _T_7334[7:0]; // @[TensorLoad.scala 259:33:@4796.4]
  assign io_tensor_rd_data_bits_6_1 = _T_7334[15:8]; // @[TensorLoad.scala 259:33:@4797.4]
  assign io_tensor_rd_data_bits_6_2 = _T_7334[23:16]; // @[TensorLoad.scala 259:33:@4798.4]
  assign io_tensor_rd_data_bits_6_3 = _T_7334[31:24]; // @[TensorLoad.scala 259:33:@4799.4]
  assign io_tensor_rd_data_bits_6_4 = _T_7334[39:32]; // @[TensorLoad.scala 259:33:@4800.4]
  assign io_tensor_rd_data_bits_6_5 = _T_7334[47:40]; // @[TensorLoad.scala 259:33:@4801.4]
  assign io_tensor_rd_data_bits_6_6 = _T_7334[55:48]; // @[TensorLoad.scala 259:33:@4802.4]
  assign io_tensor_rd_data_bits_6_7 = _T_7334[63:56]; // @[TensorLoad.scala 259:33:@4803.4]
  assign io_tensor_rd_data_bits_6_8 = _T_7334[71:64]; // @[TensorLoad.scala 259:33:@4804.4]
  assign io_tensor_rd_data_bits_6_9 = _T_7334[79:72]; // @[TensorLoad.scala 259:33:@4805.4]
  assign io_tensor_rd_data_bits_6_10 = _T_7334[87:80]; // @[TensorLoad.scala 259:33:@4806.4]
  assign io_tensor_rd_data_bits_6_11 = _T_7334[95:88]; // @[TensorLoad.scala 259:33:@4807.4]
  assign io_tensor_rd_data_bits_6_12 = _T_7334[103:96]; // @[TensorLoad.scala 259:33:@4808.4]
  assign io_tensor_rd_data_bits_6_13 = _T_7334[111:104]; // @[TensorLoad.scala 259:33:@4809.4]
  assign io_tensor_rd_data_bits_6_14 = _T_7334[119:112]; // @[TensorLoad.scala 259:33:@4810.4]
  assign io_tensor_rd_data_bits_6_15 = _T_7334[127:120]; // @[TensorLoad.scala 259:33:@4811.4]
  assign io_tensor_rd_data_bits_7_0 = _T_7476[7:0]; // @[TensorLoad.scala 259:33:@4848.4]
  assign io_tensor_rd_data_bits_7_1 = _T_7476[15:8]; // @[TensorLoad.scala 259:33:@4849.4]
  assign io_tensor_rd_data_bits_7_2 = _T_7476[23:16]; // @[TensorLoad.scala 259:33:@4850.4]
  assign io_tensor_rd_data_bits_7_3 = _T_7476[31:24]; // @[TensorLoad.scala 259:33:@4851.4]
  assign io_tensor_rd_data_bits_7_4 = _T_7476[39:32]; // @[TensorLoad.scala 259:33:@4852.4]
  assign io_tensor_rd_data_bits_7_5 = _T_7476[47:40]; // @[TensorLoad.scala 259:33:@4853.4]
  assign io_tensor_rd_data_bits_7_6 = _T_7476[55:48]; // @[TensorLoad.scala 259:33:@4854.4]
  assign io_tensor_rd_data_bits_7_7 = _T_7476[63:56]; // @[TensorLoad.scala 259:33:@4855.4]
  assign io_tensor_rd_data_bits_7_8 = _T_7476[71:64]; // @[TensorLoad.scala 259:33:@4856.4]
  assign io_tensor_rd_data_bits_7_9 = _T_7476[79:72]; // @[TensorLoad.scala 259:33:@4857.4]
  assign io_tensor_rd_data_bits_7_10 = _T_7476[87:80]; // @[TensorLoad.scala 259:33:@4858.4]
  assign io_tensor_rd_data_bits_7_11 = _T_7476[95:88]; // @[TensorLoad.scala 259:33:@4859.4]
  assign io_tensor_rd_data_bits_7_12 = _T_7476[103:96]; // @[TensorLoad.scala 259:33:@4860.4]
  assign io_tensor_rd_data_bits_7_13 = _T_7476[111:104]; // @[TensorLoad.scala 259:33:@4861.4]
  assign io_tensor_rd_data_bits_7_14 = _T_7476[119:112]; // @[TensorLoad.scala 259:33:@4862.4]
  assign io_tensor_rd_data_bits_7_15 = _T_7476[127:120]; // @[TensorLoad.scala 259:33:@4863.4]
  assign io_tensor_rd_data_bits_8_0 = _T_7618[7:0]; // @[TensorLoad.scala 259:33:@4900.4]
  assign io_tensor_rd_data_bits_8_1 = _T_7618[15:8]; // @[TensorLoad.scala 259:33:@4901.4]
  assign io_tensor_rd_data_bits_8_2 = _T_7618[23:16]; // @[TensorLoad.scala 259:33:@4902.4]
  assign io_tensor_rd_data_bits_8_3 = _T_7618[31:24]; // @[TensorLoad.scala 259:33:@4903.4]
  assign io_tensor_rd_data_bits_8_4 = _T_7618[39:32]; // @[TensorLoad.scala 259:33:@4904.4]
  assign io_tensor_rd_data_bits_8_5 = _T_7618[47:40]; // @[TensorLoad.scala 259:33:@4905.4]
  assign io_tensor_rd_data_bits_8_6 = _T_7618[55:48]; // @[TensorLoad.scala 259:33:@4906.4]
  assign io_tensor_rd_data_bits_8_7 = _T_7618[63:56]; // @[TensorLoad.scala 259:33:@4907.4]
  assign io_tensor_rd_data_bits_8_8 = _T_7618[71:64]; // @[TensorLoad.scala 259:33:@4908.4]
  assign io_tensor_rd_data_bits_8_9 = _T_7618[79:72]; // @[TensorLoad.scala 259:33:@4909.4]
  assign io_tensor_rd_data_bits_8_10 = _T_7618[87:80]; // @[TensorLoad.scala 259:33:@4910.4]
  assign io_tensor_rd_data_bits_8_11 = _T_7618[95:88]; // @[TensorLoad.scala 259:33:@4911.4]
  assign io_tensor_rd_data_bits_8_12 = _T_7618[103:96]; // @[TensorLoad.scala 259:33:@4912.4]
  assign io_tensor_rd_data_bits_8_13 = _T_7618[111:104]; // @[TensorLoad.scala 259:33:@4913.4]
  assign io_tensor_rd_data_bits_8_14 = _T_7618[119:112]; // @[TensorLoad.scala 259:33:@4914.4]
  assign io_tensor_rd_data_bits_8_15 = _T_7618[127:120]; // @[TensorLoad.scala 259:33:@4915.4]
  assign io_tensor_rd_data_bits_9_0 = _T_7760[7:0]; // @[TensorLoad.scala 259:33:@4952.4]
  assign io_tensor_rd_data_bits_9_1 = _T_7760[15:8]; // @[TensorLoad.scala 259:33:@4953.4]
  assign io_tensor_rd_data_bits_9_2 = _T_7760[23:16]; // @[TensorLoad.scala 259:33:@4954.4]
  assign io_tensor_rd_data_bits_9_3 = _T_7760[31:24]; // @[TensorLoad.scala 259:33:@4955.4]
  assign io_tensor_rd_data_bits_9_4 = _T_7760[39:32]; // @[TensorLoad.scala 259:33:@4956.4]
  assign io_tensor_rd_data_bits_9_5 = _T_7760[47:40]; // @[TensorLoad.scala 259:33:@4957.4]
  assign io_tensor_rd_data_bits_9_6 = _T_7760[55:48]; // @[TensorLoad.scala 259:33:@4958.4]
  assign io_tensor_rd_data_bits_9_7 = _T_7760[63:56]; // @[TensorLoad.scala 259:33:@4959.4]
  assign io_tensor_rd_data_bits_9_8 = _T_7760[71:64]; // @[TensorLoad.scala 259:33:@4960.4]
  assign io_tensor_rd_data_bits_9_9 = _T_7760[79:72]; // @[TensorLoad.scala 259:33:@4961.4]
  assign io_tensor_rd_data_bits_9_10 = _T_7760[87:80]; // @[TensorLoad.scala 259:33:@4962.4]
  assign io_tensor_rd_data_bits_9_11 = _T_7760[95:88]; // @[TensorLoad.scala 259:33:@4963.4]
  assign io_tensor_rd_data_bits_9_12 = _T_7760[103:96]; // @[TensorLoad.scala 259:33:@4964.4]
  assign io_tensor_rd_data_bits_9_13 = _T_7760[111:104]; // @[TensorLoad.scala 259:33:@4965.4]
  assign io_tensor_rd_data_bits_9_14 = _T_7760[119:112]; // @[TensorLoad.scala 259:33:@4966.4]
  assign io_tensor_rd_data_bits_9_15 = _T_7760[127:120]; // @[TensorLoad.scala 259:33:@4967.4]
  assign io_tensor_rd_data_bits_10_0 = _T_7902[7:0]; // @[TensorLoad.scala 259:33:@5004.4]
  assign io_tensor_rd_data_bits_10_1 = _T_7902[15:8]; // @[TensorLoad.scala 259:33:@5005.4]
  assign io_tensor_rd_data_bits_10_2 = _T_7902[23:16]; // @[TensorLoad.scala 259:33:@5006.4]
  assign io_tensor_rd_data_bits_10_3 = _T_7902[31:24]; // @[TensorLoad.scala 259:33:@5007.4]
  assign io_tensor_rd_data_bits_10_4 = _T_7902[39:32]; // @[TensorLoad.scala 259:33:@5008.4]
  assign io_tensor_rd_data_bits_10_5 = _T_7902[47:40]; // @[TensorLoad.scala 259:33:@5009.4]
  assign io_tensor_rd_data_bits_10_6 = _T_7902[55:48]; // @[TensorLoad.scala 259:33:@5010.4]
  assign io_tensor_rd_data_bits_10_7 = _T_7902[63:56]; // @[TensorLoad.scala 259:33:@5011.4]
  assign io_tensor_rd_data_bits_10_8 = _T_7902[71:64]; // @[TensorLoad.scala 259:33:@5012.4]
  assign io_tensor_rd_data_bits_10_9 = _T_7902[79:72]; // @[TensorLoad.scala 259:33:@5013.4]
  assign io_tensor_rd_data_bits_10_10 = _T_7902[87:80]; // @[TensorLoad.scala 259:33:@5014.4]
  assign io_tensor_rd_data_bits_10_11 = _T_7902[95:88]; // @[TensorLoad.scala 259:33:@5015.4]
  assign io_tensor_rd_data_bits_10_12 = _T_7902[103:96]; // @[TensorLoad.scala 259:33:@5016.4]
  assign io_tensor_rd_data_bits_10_13 = _T_7902[111:104]; // @[TensorLoad.scala 259:33:@5017.4]
  assign io_tensor_rd_data_bits_10_14 = _T_7902[119:112]; // @[TensorLoad.scala 259:33:@5018.4]
  assign io_tensor_rd_data_bits_10_15 = _T_7902[127:120]; // @[TensorLoad.scala 259:33:@5019.4]
  assign io_tensor_rd_data_bits_11_0 = _T_8044[7:0]; // @[TensorLoad.scala 259:33:@5056.4]
  assign io_tensor_rd_data_bits_11_1 = _T_8044[15:8]; // @[TensorLoad.scala 259:33:@5057.4]
  assign io_tensor_rd_data_bits_11_2 = _T_8044[23:16]; // @[TensorLoad.scala 259:33:@5058.4]
  assign io_tensor_rd_data_bits_11_3 = _T_8044[31:24]; // @[TensorLoad.scala 259:33:@5059.4]
  assign io_tensor_rd_data_bits_11_4 = _T_8044[39:32]; // @[TensorLoad.scala 259:33:@5060.4]
  assign io_tensor_rd_data_bits_11_5 = _T_8044[47:40]; // @[TensorLoad.scala 259:33:@5061.4]
  assign io_tensor_rd_data_bits_11_6 = _T_8044[55:48]; // @[TensorLoad.scala 259:33:@5062.4]
  assign io_tensor_rd_data_bits_11_7 = _T_8044[63:56]; // @[TensorLoad.scala 259:33:@5063.4]
  assign io_tensor_rd_data_bits_11_8 = _T_8044[71:64]; // @[TensorLoad.scala 259:33:@5064.4]
  assign io_tensor_rd_data_bits_11_9 = _T_8044[79:72]; // @[TensorLoad.scala 259:33:@5065.4]
  assign io_tensor_rd_data_bits_11_10 = _T_8044[87:80]; // @[TensorLoad.scala 259:33:@5066.4]
  assign io_tensor_rd_data_bits_11_11 = _T_8044[95:88]; // @[TensorLoad.scala 259:33:@5067.4]
  assign io_tensor_rd_data_bits_11_12 = _T_8044[103:96]; // @[TensorLoad.scala 259:33:@5068.4]
  assign io_tensor_rd_data_bits_11_13 = _T_8044[111:104]; // @[TensorLoad.scala 259:33:@5069.4]
  assign io_tensor_rd_data_bits_11_14 = _T_8044[119:112]; // @[TensorLoad.scala 259:33:@5070.4]
  assign io_tensor_rd_data_bits_11_15 = _T_8044[127:120]; // @[TensorLoad.scala 259:33:@5071.4]
  assign io_tensor_rd_data_bits_12_0 = _T_8186[7:0]; // @[TensorLoad.scala 259:33:@5108.4]
  assign io_tensor_rd_data_bits_12_1 = _T_8186[15:8]; // @[TensorLoad.scala 259:33:@5109.4]
  assign io_tensor_rd_data_bits_12_2 = _T_8186[23:16]; // @[TensorLoad.scala 259:33:@5110.4]
  assign io_tensor_rd_data_bits_12_3 = _T_8186[31:24]; // @[TensorLoad.scala 259:33:@5111.4]
  assign io_tensor_rd_data_bits_12_4 = _T_8186[39:32]; // @[TensorLoad.scala 259:33:@5112.4]
  assign io_tensor_rd_data_bits_12_5 = _T_8186[47:40]; // @[TensorLoad.scala 259:33:@5113.4]
  assign io_tensor_rd_data_bits_12_6 = _T_8186[55:48]; // @[TensorLoad.scala 259:33:@5114.4]
  assign io_tensor_rd_data_bits_12_7 = _T_8186[63:56]; // @[TensorLoad.scala 259:33:@5115.4]
  assign io_tensor_rd_data_bits_12_8 = _T_8186[71:64]; // @[TensorLoad.scala 259:33:@5116.4]
  assign io_tensor_rd_data_bits_12_9 = _T_8186[79:72]; // @[TensorLoad.scala 259:33:@5117.4]
  assign io_tensor_rd_data_bits_12_10 = _T_8186[87:80]; // @[TensorLoad.scala 259:33:@5118.4]
  assign io_tensor_rd_data_bits_12_11 = _T_8186[95:88]; // @[TensorLoad.scala 259:33:@5119.4]
  assign io_tensor_rd_data_bits_12_12 = _T_8186[103:96]; // @[TensorLoad.scala 259:33:@5120.4]
  assign io_tensor_rd_data_bits_12_13 = _T_8186[111:104]; // @[TensorLoad.scala 259:33:@5121.4]
  assign io_tensor_rd_data_bits_12_14 = _T_8186[119:112]; // @[TensorLoad.scala 259:33:@5122.4]
  assign io_tensor_rd_data_bits_12_15 = _T_8186[127:120]; // @[TensorLoad.scala 259:33:@5123.4]
  assign io_tensor_rd_data_bits_13_0 = _T_8328[7:0]; // @[TensorLoad.scala 259:33:@5160.4]
  assign io_tensor_rd_data_bits_13_1 = _T_8328[15:8]; // @[TensorLoad.scala 259:33:@5161.4]
  assign io_tensor_rd_data_bits_13_2 = _T_8328[23:16]; // @[TensorLoad.scala 259:33:@5162.4]
  assign io_tensor_rd_data_bits_13_3 = _T_8328[31:24]; // @[TensorLoad.scala 259:33:@5163.4]
  assign io_tensor_rd_data_bits_13_4 = _T_8328[39:32]; // @[TensorLoad.scala 259:33:@5164.4]
  assign io_tensor_rd_data_bits_13_5 = _T_8328[47:40]; // @[TensorLoad.scala 259:33:@5165.4]
  assign io_tensor_rd_data_bits_13_6 = _T_8328[55:48]; // @[TensorLoad.scala 259:33:@5166.4]
  assign io_tensor_rd_data_bits_13_7 = _T_8328[63:56]; // @[TensorLoad.scala 259:33:@5167.4]
  assign io_tensor_rd_data_bits_13_8 = _T_8328[71:64]; // @[TensorLoad.scala 259:33:@5168.4]
  assign io_tensor_rd_data_bits_13_9 = _T_8328[79:72]; // @[TensorLoad.scala 259:33:@5169.4]
  assign io_tensor_rd_data_bits_13_10 = _T_8328[87:80]; // @[TensorLoad.scala 259:33:@5170.4]
  assign io_tensor_rd_data_bits_13_11 = _T_8328[95:88]; // @[TensorLoad.scala 259:33:@5171.4]
  assign io_tensor_rd_data_bits_13_12 = _T_8328[103:96]; // @[TensorLoad.scala 259:33:@5172.4]
  assign io_tensor_rd_data_bits_13_13 = _T_8328[111:104]; // @[TensorLoad.scala 259:33:@5173.4]
  assign io_tensor_rd_data_bits_13_14 = _T_8328[119:112]; // @[TensorLoad.scala 259:33:@5174.4]
  assign io_tensor_rd_data_bits_13_15 = _T_8328[127:120]; // @[TensorLoad.scala 259:33:@5175.4]
  assign io_tensor_rd_data_bits_14_0 = _T_8470[7:0]; // @[TensorLoad.scala 259:33:@5212.4]
  assign io_tensor_rd_data_bits_14_1 = _T_8470[15:8]; // @[TensorLoad.scala 259:33:@5213.4]
  assign io_tensor_rd_data_bits_14_2 = _T_8470[23:16]; // @[TensorLoad.scala 259:33:@5214.4]
  assign io_tensor_rd_data_bits_14_3 = _T_8470[31:24]; // @[TensorLoad.scala 259:33:@5215.4]
  assign io_tensor_rd_data_bits_14_4 = _T_8470[39:32]; // @[TensorLoad.scala 259:33:@5216.4]
  assign io_tensor_rd_data_bits_14_5 = _T_8470[47:40]; // @[TensorLoad.scala 259:33:@5217.4]
  assign io_tensor_rd_data_bits_14_6 = _T_8470[55:48]; // @[TensorLoad.scala 259:33:@5218.4]
  assign io_tensor_rd_data_bits_14_7 = _T_8470[63:56]; // @[TensorLoad.scala 259:33:@5219.4]
  assign io_tensor_rd_data_bits_14_8 = _T_8470[71:64]; // @[TensorLoad.scala 259:33:@5220.4]
  assign io_tensor_rd_data_bits_14_9 = _T_8470[79:72]; // @[TensorLoad.scala 259:33:@5221.4]
  assign io_tensor_rd_data_bits_14_10 = _T_8470[87:80]; // @[TensorLoad.scala 259:33:@5222.4]
  assign io_tensor_rd_data_bits_14_11 = _T_8470[95:88]; // @[TensorLoad.scala 259:33:@5223.4]
  assign io_tensor_rd_data_bits_14_12 = _T_8470[103:96]; // @[TensorLoad.scala 259:33:@5224.4]
  assign io_tensor_rd_data_bits_14_13 = _T_8470[111:104]; // @[TensorLoad.scala 259:33:@5225.4]
  assign io_tensor_rd_data_bits_14_14 = _T_8470[119:112]; // @[TensorLoad.scala 259:33:@5226.4]
  assign io_tensor_rd_data_bits_14_15 = _T_8470[127:120]; // @[TensorLoad.scala 259:33:@5227.4]
  assign io_tensor_rd_data_bits_15_0 = _T_8612[7:0]; // @[TensorLoad.scala 259:33:@5264.4]
  assign io_tensor_rd_data_bits_15_1 = _T_8612[15:8]; // @[TensorLoad.scala 259:33:@5265.4]
  assign io_tensor_rd_data_bits_15_2 = _T_8612[23:16]; // @[TensorLoad.scala 259:33:@5266.4]
  assign io_tensor_rd_data_bits_15_3 = _T_8612[31:24]; // @[TensorLoad.scala 259:33:@5267.4]
  assign io_tensor_rd_data_bits_15_4 = _T_8612[39:32]; // @[TensorLoad.scala 259:33:@5268.4]
  assign io_tensor_rd_data_bits_15_5 = _T_8612[47:40]; // @[TensorLoad.scala 259:33:@5269.4]
  assign io_tensor_rd_data_bits_15_6 = _T_8612[55:48]; // @[TensorLoad.scala 259:33:@5270.4]
  assign io_tensor_rd_data_bits_15_7 = _T_8612[63:56]; // @[TensorLoad.scala 259:33:@5271.4]
  assign io_tensor_rd_data_bits_15_8 = _T_8612[71:64]; // @[TensorLoad.scala 259:33:@5272.4]
  assign io_tensor_rd_data_bits_15_9 = _T_8612[79:72]; // @[TensorLoad.scala 259:33:@5273.4]
  assign io_tensor_rd_data_bits_15_10 = _T_8612[87:80]; // @[TensorLoad.scala 259:33:@5274.4]
  assign io_tensor_rd_data_bits_15_11 = _T_8612[95:88]; // @[TensorLoad.scala 259:33:@5275.4]
  assign io_tensor_rd_data_bits_15_12 = _T_8612[103:96]; // @[TensorLoad.scala 259:33:@5276.4]
  assign io_tensor_rd_data_bits_15_13 = _T_8612[111:104]; // @[TensorLoad.scala 259:33:@5277.4]
  assign io_tensor_rd_data_bits_15_14 = _T_8612[119:112]; // @[TensorLoad.scala 259:33:@5278.4]
  assign io_tensor_rd_data_bits_15_15 = _T_8612[127:120]; // @[TensorLoad.scala 259:33:@5279.4]
  assign dataCtrl_clock = clock; // @[:@3168.4]
  assign dataCtrl_io_start = _T_4420 & io_start; // @[TensorLoad.scala 147:21:@3303.4]
  assign dataCtrl_io_inst = io_inst; // @[TensorLoad.scala 148:20:@3304.4]
  assign dataCtrl_io_baddr = io_baddr; // @[TensorLoad.scala 149:21:@3305.4]
  assign dataCtrl_io_xinit = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[TensorLoad.scala 150:21:@3307.4]
  assign dataCtrl_io_xupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 151:23:@3309.4]
  assign dataCtrl_io_yupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 152:23:@3311.4]
  assign yPadCtrl0_clock = clock; // @[:@3172.4]
  assign yPadCtrl0_reset = reset; // @[:@3173.4]
  assign yPadCtrl0_io_start = _T_4433 & io_start; // @[TensorLoad.scala 161:22:@3326.4]
  assign yPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 176:21:@3368.4]
  assign yPadCtrl1_clock = clock; // @[:@3175.4]
  assign yPadCtrl1_reset = reset; // @[:@3176.4]
  assign yPadCtrl1_io_start = _T_4408 & _T_4445; // @[TensorLoad.scala 163:22:@3337.4]
  assign yPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 177:21:@3369.4]
  assign xPadCtrl0_clock = clock; // @[:@3178.4]
  assign xPadCtrl0_reset = reset; // @[:@3179.4]
  assign xPadCtrl0_io_start = _T_4398 & _T_4466; // @[TensorLoad.scala 167:22:@3357.4]
  assign xPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 178:21:@3370.4]
  assign xPadCtrl1_clock = clock; // @[:@3181.4]
  assign xPadCtrl1_reset = reset; // @[:@3182.4]
  assign xPadCtrl1_io_start = _T_4471 & _T_4477; // @[TensorLoad.scala 173:22:@3367.4]
  assign xPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 179:21:@3371.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_0_0[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_0_1[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_1_0[initvar] = _RAND_2[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_1_1[initvar] = _RAND_3[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_2_0[initvar] = _RAND_4[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_2_1[initvar] = _RAND_5[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_3_0[initvar] = _RAND_6[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_3_1[initvar] = _RAND_7[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_4_0[initvar] = _RAND_8[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_4_1[initvar] = _RAND_9[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_5_0[initvar] = _RAND_10[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_5_1[initvar] = _RAND_11[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_12 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_6_0[initvar] = _RAND_12[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_6_1[initvar] = _RAND_13[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_14 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_7_0[initvar] = _RAND_14[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_15 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_7_1[initvar] = _RAND_15[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_16 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_8_0[initvar] = _RAND_16[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_8_1[initvar] = _RAND_17[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_18 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_9_0[initvar] = _RAND_18[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_19 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_9_1[initvar] = _RAND_19[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_20 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_10_0[initvar] = _RAND_20[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_10_1[initvar] = _RAND_21[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_22 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_11_0[initvar] = _RAND_22[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_23 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_11_1[initvar] = _RAND_23[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_24 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_12_0[initvar] = _RAND_24[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_12_1[initvar] = _RAND_25[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_26 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_13_0[initvar] = _RAND_26[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_27 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_13_1[initvar] = _RAND_27[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_28 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_14_0[initvar] = _RAND_28[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_14_1[initvar] = _RAND_29[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_30 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_15_0[initvar] = _RAND_30[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_31 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_15_1[initvar] = _RAND_31[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  dataCtrlDone = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  tag = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  set = _RAND_34[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  state = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  waddr_cur = _RAND_36[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  waddr_nxt = _RAND_37[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  rvalid = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  tensorFile_0_0_rdata_0_addr_pipe_0 = _RAND_39[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  tensorFile_0_1_rdata_0_addr_pipe_0 = _RAND_40[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  tensorFile_1_0_rdata_1_addr_pipe_0 = _RAND_41[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  tensorFile_1_1_rdata_1_addr_pipe_0 = _RAND_42[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  tensorFile_2_0_rdata_2_addr_pipe_0 = _RAND_43[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  tensorFile_2_1_rdata_2_addr_pipe_0 = _RAND_44[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  tensorFile_3_0_rdata_3_addr_pipe_0 = _RAND_45[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  tensorFile_3_1_rdata_3_addr_pipe_0 = _RAND_46[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  tensorFile_4_0_rdata_4_addr_pipe_0 = _RAND_47[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  tensorFile_4_1_rdata_4_addr_pipe_0 = _RAND_48[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  tensorFile_5_0_rdata_5_addr_pipe_0 = _RAND_49[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  tensorFile_5_1_rdata_5_addr_pipe_0 = _RAND_50[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  tensorFile_6_0_rdata_6_addr_pipe_0 = _RAND_51[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  tensorFile_6_1_rdata_6_addr_pipe_0 = _RAND_52[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  tensorFile_7_0_rdata_7_addr_pipe_0 = _RAND_53[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  tensorFile_7_1_rdata_7_addr_pipe_0 = _RAND_54[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  tensorFile_8_0_rdata_8_addr_pipe_0 = _RAND_55[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  tensorFile_8_1_rdata_8_addr_pipe_0 = _RAND_56[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  tensorFile_9_0_rdata_9_addr_pipe_0 = _RAND_57[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  tensorFile_9_1_rdata_9_addr_pipe_0 = _RAND_58[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  tensorFile_10_0_rdata_10_addr_pipe_0 = _RAND_59[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  tensorFile_10_1_rdata_10_addr_pipe_0 = _RAND_60[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  tensorFile_11_0_rdata_11_addr_pipe_0 = _RAND_61[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  tensorFile_11_1_rdata_11_addr_pipe_0 = _RAND_62[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  tensorFile_12_0_rdata_12_addr_pipe_0 = _RAND_63[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  tensorFile_12_1_rdata_12_addr_pipe_0 = _RAND_64[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  tensorFile_13_0_rdata_13_addr_pipe_0 = _RAND_65[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  tensorFile_13_1_rdata_13_addr_pipe_0 = _RAND_66[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  tensorFile_14_0_rdata_14_addr_pipe_0 = _RAND_67[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  tensorFile_14_1_rdata_14_addr_pipe_0 = _RAND_68[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  tensorFile_15_0_rdata_15_addr_pipe_0 = _RAND_69[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  tensorFile_15_1_rdata_15_addr_pipe_0 = _RAND_70[9:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tensorFile_0_0__T_4976_en & tensorFile_0_0__T_4976_mask) begin
      tensorFile_0_0[tensorFile_0_0__T_4976_addr] <= tensorFile_0_0__T_4976_data; // @[TensorLoad.scala 222:16:@3450.4]
    end
    if(tensorFile_0_1__T_4976_en & tensorFile_0_1__T_4976_mask) begin
      tensorFile_0_1[tensorFile_0_1__T_4976_addr] <= tensorFile_0_1__T_4976_data; // @[TensorLoad.scala 222:16:@3450.4]
    end
    if(tensorFile_1_0__T_5063_en & tensorFile_1_0__T_5063_mask) begin
      tensorFile_1_0[tensorFile_1_0__T_5063_addr] <= tensorFile_1_0__T_5063_data; // @[TensorLoad.scala 222:16:@3451.4]
    end
    if(tensorFile_1_1__T_5063_en & tensorFile_1_1__T_5063_mask) begin
      tensorFile_1_1[tensorFile_1_1__T_5063_addr] <= tensorFile_1_1__T_5063_data; // @[TensorLoad.scala 222:16:@3451.4]
    end
    if(tensorFile_2_0__T_5150_en & tensorFile_2_0__T_5150_mask) begin
      tensorFile_2_0[tensorFile_2_0__T_5150_addr] <= tensorFile_2_0__T_5150_data; // @[TensorLoad.scala 222:16:@3452.4]
    end
    if(tensorFile_2_1__T_5150_en & tensorFile_2_1__T_5150_mask) begin
      tensorFile_2_1[tensorFile_2_1__T_5150_addr] <= tensorFile_2_1__T_5150_data; // @[TensorLoad.scala 222:16:@3452.4]
    end
    if(tensorFile_3_0__T_5237_en & tensorFile_3_0__T_5237_mask) begin
      tensorFile_3_0[tensorFile_3_0__T_5237_addr] <= tensorFile_3_0__T_5237_data; // @[TensorLoad.scala 222:16:@3453.4]
    end
    if(tensorFile_3_1__T_5237_en & tensorFile_3_1__T_5237_mask) begin
      tensorFile_3_1[tensorFile_3_1__T_5237_addr] <= tensorFile_3_1__T_5237_data; // @[TensorLoad.scala 222:16:@3453.4]
    end
    if(tensorFile_4_0__T_5324_en & tensorFile_4_0__T_5324_mask) begin
      tensorFile_4_0[tensorFile_4_0__T_5324_addr] <= tensorFile_4_0__T_5324_data; // @[TensorLoad.scala 222:16:@3454.4]
    end
    if(tensorFile_4_1__T_5324_en & tensorFile_4_1__T_5324_mask) begin
      tensorFile_4_1[tensorFile_4_1__T_5324_addr] <= tensorFile_4_1__T_5324_data; // @[TensorLoad.scala 222:16:@3454.4]
    end
    if(tensorFile_5_0__T_5411_en & tensorFile_5_0__T_5411_mask) begin
      tensorFile_5_0[tensorFile_5_0__T_5411_addr] <= tensorFile_5_0__T_5411_data; // @[TensorLoad.scala 222:16:@3455.4]
    end
    if(tensorFile_5_1__T_5411_en & tensorFile_5_1__T_5411_mask) begin
      tensorFile_5_1[tensorFile_5_1__T_5411_addr] <= tensorFile_5_1__T_5411_data; // @[TensorLoad.scala 222:16:@3455.4]
    end
    if(tensorFile_6_0__T_5498_en & tensorFile_6_0__T_5498_mask) begin
      tensorFile_6_0[tensorFile_6_0__T_5498_addr] <= tensorFile_6_0__T_5498_data; // @[TensorLoad.scala 222:16:@3456.4]
    end
    if(tensorFile_6_1__T_5498_en & tensorFile_6_1__T_5498_mask) begin
      tensorFile_6_1[tensorFile_6_1__T_5498_addr] <= tensorFile_6_1__T_5498_data; // @[TensorLoad.scala 222:16:@3456.4]
    end
    if(tensorFile_7_0__T_5585_en & tensorFile_7_0__T_5585_mask) begin
      tensorFile_7_0[tensorFile_7_0__T_5585_addr] <= tensorFile_7_0__T_5585_data; // @[TensorLoad.scala 222:16:@3457.4]
    end
    if(tensorFile_7_1__T_5585_en & tensorFile_7_1__T_5585_mask) begin
      tensorFile_7_1[tensorFile_7_1__T_5585_addr] <= tensorFile_7_1__T_5585_data; // @[TensorLoad.scala 222:16:@3457.4]
    end
    if(tensorFile_8_0__T_5672_en & tensorFile_8_0__T_5672_mask) begin
      tensorFile_8_0[tensorFile_8_0__T_5672_addr] <= tensorFile_8_0__T_5672_data; // @[TensorLoad.scala 222:16:@3458.4]
    end
    if(tensorFile_8_1__T_5672_en & tensorFile_8_1__T_5672_mask) begin
      tensorFile_8_1[tensorFile_8_1__T_5672_addr] <= tensorFile_8_1__T_5672_data; // @[TensorLoad.scala 222:16:@3458.4]
    end
    if(tensorFile_9_0__T_5759_en & tensorFile_9_0__T_5759_mask) begin
      tensorFile_9_0[tensorFile_9_0__T_5759_addr] <= tensorFile_9_0__T_5759_data; // @[TensorLoad.scala 222:16:@3459.4]
    end
    if(tensorFile_9_1__T_5759_en & tensorFile_9_1__T_5759_mask) begin
      tensorFile_9_1[tensorFile_9_1__T_5759_addr] <= tensorFile_9_1__T_5759_data; // @[TensorLoad.scala 222:16:@3459.4]
    end
    if(tensorFile_10_0__T_5846_en & tensorFile_10_0__T_5846_mask) begin
      tensorFile_10_0[tensorFile_10_0__T_5846_addr] <= tensorFile_10_0__T_5846_data; // @[TensorLoad.scala 222:16:@3460.4]
    end
    if(tensorFile_10_1__T_5846_en & tensorFile_10_1__T_5846_mask) begin
      tensorFile_10_1[tensorFile_10_1__T_5846_addr] <= tensorFile_10_1__T_5846_data; // @[TensorLoad.scala 222:16:@3460.4]
    end
    if(tensorFile_11_0__T_5933_en & tensorFile_11_0__T_5933_mask) begin
      tensorFile_11_0[tensorFile_11_0__T_5933_addr] <= tensorFile_11_0__T_5933_data; // @[TensorLoad.scala 222:16:@3461.4]
    end
    if(tensorFile_11_1__T_5933_en & tensorFile_11_1__T_5933_mask) begin
      tensorFile_11_1[tensorFile_11_1__T_5933_addr] <= tensorFile_11_1__T_5933_data; // @[TensorLoad.scala 222:16:@3461.4]
    end
    if(tensorFile_12_0__T_6020_en & tensorFile_12_0__T_6020_mask) begin
      tensorFile_12_0[tensorFile_12_0__T_6020_addr] <= tensorFile_12_0__T_6020_data; // @[TensorLoad.scala 222:16:@3462.4]
    end
    if(tensorFile_12_1__T_6020_en & tensorFile_12_1__T_6020_mask) begin
      tensorFile_12_1[tensorFile_12_1__T_6020_addr] <= tensorFile_12_1__T_6020_data; // @[TensorLoad.scala 222:16:@3462.4]
    end
    if(tensorFile_13_0__T_6107_en & tensorFile_13_0__T_6107_mask) begin
      tensorFile_13_0[tensorFile_13_0__T_6107_addr] <= tensorFile_13_0__T_6107_data; // @[TensorLoad.scala 222:16:@3463.4]
    end
    if(tensorFile_13_1__T_6107_en & tensorFile_13_1__T_6107_mask) begin
      tensorFile_13_1[tensorFile_13_1__T_6107_addr] <= tensorFile_13_1__T_6107_data; // @[TensorLoad.scala 222:16:@3463.4]
    end
    if(tensorFile_14_0__T_6194_en & tensorFile_14_0__T_6194_mask) begin
      tensorFile_14_0[tensorFile_14_0__T_6194_addr] <= tensorFile_14_0__T_6194_data; // @[TensorLoad.scala 222:16:@3464.4]
    end
    if(tensorFile_14_1__T_6194_en & tensorFile_14_1__T_6194_mask) begin
      tensorFile_14_1[tensorFile_14_1__T_6194_addr] <= tensorFile_14_1__T_6194_data; // @[TensorLoad.scala 222:16:@3464.4]
    end
    if(tensorFile_15_0__T_6281_en & tensorFile_15_0__T_6281_mask) begin
      tensorFile_15_0[tensorFile_15_0__T_6281_addr] <= tensorFile_15_0__T_6281_data; // @[TensorLoad.scala 222:16:@3465.4]
    end
    if(tensorFile_15_1__T_6281_en & tensorFile_15_1__T_6281_mask) begin
      tensorFile_15_1[tensorFile_15_1__T_6281_addr] <= tensorFile_15_1__T_6281_data; // @[TensorLoad.scala 222:16:@3465.4]
    end
    if (reset) begin
      dataCtrlDone <= 1'h0;
    end else begin
      if (_T_4420) begin
        dataCtrlDone <= 1'h0;
      end else begin
        if (_T_4428) begin
          dataCtrlDone <= 1'h1;
        end
      end
    end
    if (_T_4492) begin
      tag <= 1'h0;
    end else begin
      if (_T_4495) begin
        tag <= _T_4498;
      end
    end
    if (_T_4506) begin
      set <= 4'h0;
    end else begin
      if (_T_4512) begin
        set <= _T_4515;
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_4394) begin
        if (io_start) begin
          if (_T_4396) begin
            state <= 3'h1;
          end else begin
            if (_T_4398) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end
      end else begin
        if (_T_4399) begin
          if (yPadCtrl0_io_done) begin
            if (_T_4398) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end else begin
          if (_T_4402) begin
            if (xPadCtrl0_io_done) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_4403) begin
              if (io_vme_rd_cmd_ready) begin
                state <= 3'h4;
              end
            end else begin
              if (_T_4404) begin
                if (io_vme_rd_data_valid) begin
                  if (dataCtrl_io_done) begin
                    if (_T_4406) begin
                      state <= 3'h5;
                    end else begin
                      if (_T_4408) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end
                  end else begin
                    if (dataCtrl_io_stride) begin
                      if (_T_4406) begin
                        state <= 3'h5;
                      end else begin
                        if (_T_4398) begin
                          state <= 3'h2;
                        end else begin
                          state <= 3'h3;
                        end
                      end
                    end else begin
                      if (dataCtrl_io_split) begin
                        state <= 3'h3;
                      end
                    end
                  end
                end
              end else begin
                if (_T_4413) begin
                  if (xPadCtrl1_io_done) begin
                    if (dataCtrlDone) begin
                      if (_T_4408) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end else begin
                      if (_T_4398) begin
                        state <= 3'h2;
                      end else begin
                        state <= 3'h3;
                      end
                    end
                  end
                end else begin
                  if (_T_4418) begin
                    if (_T_4419) begin
                      state <= 3'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    waddr_cur <= _GEN_37[9:0];
    waddr_nxt <= _GEN_38[9:0];
    rvalid <= io_tensor_rd_idx_valid;
    if (_GEN_216) begin
      tensorFile_0_0_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_0_1_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_1_0_rdata_1_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_1_1_rdata_1_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_2_0_rdata_2_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_2_1_rdata_2_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_3_0_rdata_3_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_3_1_rdata_3_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_4_0_rdata_4_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_4_1_rdata_4_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_5_0_rdata_5_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_5_1_rdata_5_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_6_0_rdata_6_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_6_1_rdata_6_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_7_0_rdata_7_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_7_1_rdata_7_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_8_0_rdata_8_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_8_1_rdata_8_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_9_0_rdata_9_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_9_1_rdata_9_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_10_0_rdata_10_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_10_1_rdata_10_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_11_0_rdata_11_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_11_1_rdata_11_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_12_0_rdata_12_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_12_1_rdata_12_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_13_0_rdata_13_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_13_1_rdata_13_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_14_0_rdata_14_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_14_1_rdata_14_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_15_0_rdata_15_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_216) begin
      tensorFile_15_1_rdata_15_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
  end
endmodule
module Load( // @[:@5298.2]
  input          clock, // @[:@5299.4]
  input          reset, // @[:@5300.4]
  input          io_i_post, // @[:@5301.4]
  output         io_o_post, // @[:@5301.4]
  output         io_inst_ready, // @[:@5301.4]
  input          io_inst_valid, // @[:@5301.4]
  input  [127:0] io_inst_bits, // @[:@5301.4]
  input  [31:0]  io_inp_baddr, // @[:@5301.4]
  input  [31:0]  io_wgt_baddr, // @[:@5301.4]
  input          io_vme_rd_0_cmd_ready, // @[:@5301.4]
  output         io_vme_rd_0_cmd_valid, // @[:@5301.4]
  output [31:0]  io_vme_rd_0_cmd_bits_addr, // @[:@5301.4]
  output [7:0]   io_vme_rd_0_cmd_bits_len, // @[:@5301.4]
  output         io_vme_rd_0_data_ready, // @[:@5301.4]
  input          io_vme_rd_0_data_valid, // @[:@5301.4]
  input  [63:0]  io_vme_rd_0_data_bits, // @[:@5301.4]
  input          io_vme_rd_1_cmd_ready, // @[:@5301.4]
  output         io_vme_rd_1_cmd_valid, // @[:@5301.4]
  output [31:0]  io_vme_rd_1_cmd_bits_addr, // @[:@5301.4]
  output [7:0]   io_vme_rd_1_cmd_bits_len, // @[:@5301.4]
  output         io_vme_rd_1_data_ready, // @[:@5301.4]
  input          io_vme_rd_1_data_valid, // @[:@5301.4]
  input  [63:0]  io_vme_rd_1_data_bits, // @[:@5301.4]
  input          io_inp_rd_idx_valid, // @[:@5301.4]
  input  [10:0]  io_inp_rd_idx_bits, // @[:@5301.4]
  output         io_inp_rd_data_valid, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_0, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_1, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_2, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_3, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_4, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_5, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_6, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_7, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_8, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_9, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_10, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_11, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_12, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_13, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_14, // @[:@5301.4]
  output [7:0]   io_inp_rd_data_bits_0_15, // @[:@5301.4]
  input          io_wgt_rd_idx_valid, // @[:@5301.4]
  input  [9:0]   io_wgt_rd_idx_bits, // @[:@5301.4]
  output         io_wgt_rd_data_valid, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_0_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_1_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_2_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_3_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_4_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_5_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_6_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_7_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_8_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_9_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_10_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_11_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_12_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_13_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_14_15, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_0, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_1, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_2, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_3, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_4, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_5, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_6, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_7, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_8, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_9, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_10, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_11, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_12, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_13, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_14, // @[:@5301.4]
  output [7:0]   io_wgt_rd_data_bits_15_15 // @[:@5301.4]
);
  wire  s_clock; // @[Load.scala 49:17:@5304.4]
  wire  s_reset; // @[Load.scala 49:17:@5304.4]
  wire  s_io_spost; // @[Load.scala 49:17:@5304.4]
  wire  s_io_swait; // @[Load.scala 49:17:@5304.4]
  wire  s_io_sready; // @[Load.scala 49:17:@5304.4]
  wire  inst_q_clock; // @[Load.scala 50:22:@5307.4]
  wire  inst_q_reset; // @[Load.scala 50:22:@5307.4]
  wire  inst_q_io_enq_ready; // @[Load.scala 50:22:@5307.4]
  wire  inst_q_io_enq_valid; // @[Load.scala 50:22:@5307.4]
  wire [127:0] inst_q_io_enq_bits; // @[Load.scala 50:22:@5307.4]
  wire  inst_q_io_deq_ready; // @[Load.scala 50:22:@5307.4]
  wire  inst_q_io_deq_valid; // @[Load.scala 50:22:@5307.4]
  wire [127:0] inst_q_io_deq_bits; // @[Load.scala 50:22:@5307.4]
  wire [127:0] dec_io_inst; // @[Load.scala 52:19:@5310.4]
  wire  dec_io_push_next; // @[Load.scala 52:19:@5310.4]
  wire  dec_io_pop_next; // @[Load.scala 52:19:@5310.4]
  wire  dec_io_isInput; // @[Load.scala 52:19:@5310.4]
  wire  dec_io_isWeight; // @[Load.scala 52:19:@5310.4]
  wire  dec_io_isSync; // @[Load.scala 52:19:@5310.4]
  wire  tensorLoad_0_clock; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_0_reset; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_0_io_start; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_0_io_done; // @[Load.scala 58:32:@5314.4]
  wire [127:0] tensorLoad_0_io_inst; // @[Load.scala 58:32:@5314.4]
  wire [31:0] tensorLoad_0_io_baddr; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_0_io_vme_rd_cmd_ready; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_0_io_vme_rd_cmd_valid; // @[Load.scala 58:32:@5314.4]
  wire [31:0] tensorLoad_0_io_vme_rd_cmd_bits_addr; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_vme_rd_cmd_bits_len; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_0_io_vme_rd_data_ready; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_0_io_vme_rd_data_valid; // @[Load.scala 58:32:@5314.4]
  wire [63:0] tensorLoad_0_io_vme_rd_data_bits; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_0_io_tensor_rd_idx_valid; // @[Load.scala 58:32:@5314.4]
  wire [10:0] tensorLoad_0_io_tensor_rd_idx_bits; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_0_io_tensor_rd_data_valid; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_0; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_1; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_2; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_3; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_4; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_5; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_6; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_7; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_8; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_9; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_10; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_11; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_12; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_13; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_14; // @[Load.scala 58:32:@5314.4]
  wire [7:0] tensorLoad_0_io_tensor_rd_data_bits_0_15; // @[Load.scala 58:32:@5314.4]
  wire  tensorLoad_1_clock; // @[Load.scala 58:32:@5317.4]
  wire  tensorLoad_1_reset; // @[Load.scala 58:32:@5317.4]
  wire  tensorLoad_1_io_start; // @[Load.scala 58:32:@5317.4]
  wire  tensorLoad_1_io_done; // @[Load.scala 58:32:@5317.4]
  wire [127:0] tensorLoad_1_io_inst; // @[Load.scala 58:32:@5317.4]
  wire [31:0] tensorLoad_1_io_baddr; // @[Load.scala 58:32:@5317.4]
  wire  tensorLoad_1_io_vme_rd_cmd_ready; // @[Load.scala 58:32:@5317.4]
  wire  tensorLoad_1_io_vme_rd_cmd_valid; // @[Load.scala 58:32:@5317.4]
  wire [31:0] tensorLoad_1_io_vme_rd_cmd_bits_addr; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_vme_rd_cmd_bits_len; // @[Load.scala 58:32:@5317.4]
  wire  tensorLoad_1_io_vme_rd_data_ready; // @[Load.scala 58:32:@5317.4]
  wire  tensorLoad_1_io_vme_rd_data_valid; // @[Load.scala 58:32:@5317.4]
  wire [63:0] tensorLoad_1_io_vme_rd_data_bits; // @[Load.scala 58:32:@5317.4]
  wire  tensorLoad_1_io_tensor_rd_idx_valid; // @[Load.scala 58:32:@5317.4]
  wire [9:0] tensorLoad_1_io_tensor_rd_idx_bits; // @[Load.scala 58:32:@5317.4]
  wire  tensorLoad_1_io_tensor_rd_data_valid; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_0_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_1_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_2_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_3_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_4_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_5_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_6_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_7_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_8_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_9_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_10_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_11_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_12_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_13_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_14_15; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_0; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_1; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_2; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_3; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_4; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_5; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_6; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_7; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_8; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_9; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_10; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_11; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_12; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_13; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_14; // @[Load.scala 58:32:@5317.4]
  wire [7:0] tensorLoad_1_io_tensor_rd_data_bits_15_15; // @[Load.scala 58:32:@5317.4]
  reg [1:0] state; // @[Load.scala 47:22:@5303.4]
  reg [31:0] _RAND_0;
  wire  _T_4999; // @[Load.scala 60:40:@5320.4]
  wire  start; // @[Load.scala 60:35:@5321.4]
  wire  done; // @[Load.scala 61:17:@5322.4]
  wire  _T_5000; // @[Conditional.scala 37:30:@5323.4]
  wire  _T_5001; // @[Load.scala 69:35:@5330.10]
  wire [1:0] _GEN_0; // @[Load.scala 69:55:@5331.10]
  wire [1:0] _GEN_1; // @[Load.scala 67:29:@5326.8]
  wire [1:0] _GEN_2; // @[Load.scala 66:19:@5325.6]
  wire  _T_5002; // @[Conditional.scala 37:30:@5337.6]
  wire  _T_5003; // @[Conditional.scala 37:30:@5342.8]
  wire [1:0] _GEN_3; // @[Load.scala 78:18:@5344.10]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@5343.8]
  wire [1:0] _GEN_5; // @[Conditional.scala 39:67:@5338.6]
  wire [1:0] _GEN_6; // @[Conditional.scala 40:58:@5324.4]
  wire  _T_5004; // @[Load.scala 86:33:@5351.4]
  wire  _T_5005; // @[Load.scala 86:42:@5352.4]
  wire  _T_5006; // @[Load.scala 86:59:@5353.4]
  wire  _T_5007; // @[Load.scala 86:50:@5354.4]
  wire  _T_5008; // @[Load.scala 94:37:@5356.4]
  wire  _T_5009; // @[Load.scala 94:47:@5357.4]
  Semaphore s ( // @[Load.scala 49:17:@5304.4]
    .clock(s_clock),
    .reset(s_reset),
    .io_spost(s_io_spost),
    .io_swait(s_io_swait),
    .io_sready(s_io_sready)
  );
  Queue_1 inst_q ( // @[Load.scala 50:22:@5307.4]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits)
  );
  LoadDecode dec ( // @[Load.scala 52:19:@5310.4]
    .io_inst(dec_io_inst),
    .io_push_next(dec_io_push_next),
    .io_pop_next(dec_io_pop_next),
    .io_isInput(dec_io_isInput),
    .io_isWeight(dec_io_isWeight),
    .io_isSync(dec_io_isSync)
  );
  TensorLoad tensorLoad_0 ( // @[Load.scala 58:32:@5314.4]
    .clock(tensorLoad_0_clock),
    .reset(tensorLoad_0_reset),
    .io_start(tensorLoad_0_io_start),
    .io_done(tensorLoad_0_io_done),
    .io_inst(tensorLoad_0_io_inst),
    .io_baddr(tensorLoad_0_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_0_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_0_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_0_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_0_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(tensorLoad_0_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorLoad_0_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(tensorLoad_0_io_vme_rd_data_bits),
    .io_tensor_rd_idx_valid(tensorLoad_0_io_tensor_rd_idx_valid),
    .io_tensor_rd_idx_bits(tensorLoad_0_io_tensor_rd_idx_bits),
    .io_tensor_rd_data_valid(tensorLoad_0_io_tensor_rd_data_valid),
    .io_tensor_rd_data_bits_0_0(tensorLoad_0_io_tensor_rd_data_bits_0_0),
    .io_tensor_rd_data_bits_0_1(tensorLoad_0_io_tensor_rd_data_bits_0_1),
    .io_tensor_rd_data_bits_0_2(tensorLoad_0_io_tensor_rd_data_bits_0_2),
    .io_tensor_rd_data_bits_0_3(tensorLoad_0_io_tensor_rd_data_bits_0_3),
    .io_tensor_rd_data_bits_0_4(tensorLoad_0_io_tensor_rd_data_bits_0_4),
    .io_tensor_rd_data_bits_0_5(tensorLoad_0_io_tensor_rd_data_bits_0_5),
    .io_tensor_rd_data_bits_0_6(tensorLoad_0_io_tensor_rd_data_bits_0_6),
    .io_tensor_rd_data_bits_0_7(tensorLoad_0_io_tensor_rd_data_bits_0_7),
    .io_tensor_rd_data_bits_0_8(tensorLoad_0_io_tensor_rd_data_bits_0_8),
    .io_tensor_rd_data_bits_0_9(tensorLoad_0_io_tensor_rd_data_bits_0_9),
    .io_tensor_rd_data_bits_0_10(tensorLoad_0_io_tensor_rd_data_bits_0_10),
    .io_tensor_rd_data_bits_0_11(tensorLoad_0_io_tensor_rd_data_bits_0_11),
    .io_tensor_rd_data_bits_0_12(tensorLoad_0_io_tensor_rd_data_bits_0_12),
    .io_tensor_rd_data_bits_0_13(tensorLoad_0_io_tensor_rd_data_bits_0_13),
    .io_tensor_rd_data_bits_0_14(tensorLoad_0_io_tensor_rd_data_bits_0_14),
    .io_tensor_rd_data_bits_0_15(tensorLoad_0_io_tensor_rd_data_bits_0_15)
  );
  TensorLoad_1 tensorLoad_1 ( // @[Load.scala 58:32:@5317.4]
    .clock(tensorLoad_1_clock),
    .reset(tensorLoad_1_reset),
    .io_start(tensorLoad_1_io_start),
    .io_done(tensorLoad_1_io_done),
    .io_inst(tensorLoad_1_io_inst),
    .io_baddr(tensorLoad_1_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_1_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_1_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_1_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_1_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(tensorLoad_1_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorLoad_1_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(tensorLoad_1_io_vme_rd_data_bits),
    .io_tensor_rd_idx_valid(tensorLoad_1_io_tensor_rd_idx_valid),
    .io_tensor_rd_idx_bits(tensorLoad_1_io_tensor_rd_idx_bits),
    .io_tensor_rd_data_valid(tensorLoad_1_io_tensor_rd_data_valid),
    .io_tensor_rd_data_bits_0_0(tensorLoad_1_io_tensor_rd_data_bits_0_0),
    .io_tensor_rd_data_bits_0_1(tensorLoad_1_io_tensor_rd_data_bits_0_1),
    .io_tensor_rd_data_bits_0_2(tensorLoad_1_io_tensor_rd_data_bits_0_2),
    .io_tensor_rd_data_bits_0_3(tensorLoad_1_io_tensor_rd_data_bits_0_3),
    .io_tensor_rd_data_bits_0_4(tensorLoad_1_io_tensor_rd_data_bits_0_4),
    .io_tensor_rd_data_bits_0_5(tensorLoad_1_io_tensor_rd_data_bits_0_5),
    .io_tensor_rd_data_bits_0_6(tensorLoad_1_io_tensor_rd_data_bits_0_6),
    .io_tensor_rd_data_bits_0_7(tensorLoad_1_io_tensor_rd_data_bits_0_7),
    .io_tensor_rd_data_bits_0_8(tensorLoad_1_io_tensor_rd_data_bits_0_8),
    .io_tensor_rd_data_bits_0_9(tensorLoad_1_io_tensor_rd_data_bits_0_9),
    .io_tensor_rd_data_bits_0_10(tensorLoad_1_io_tensor_rd_data_bits_0_10),
    .io_tensor_rd_data_bits_0_11(tensorLoad_1_io_tensor_rd_data_bits_0_11),
    .io_tensor_rd_data_bits_0_12(tensorLoad_1_io_tensor_rd_data_bits_0_12),
    .io_tensor_rd_data_bits_0_13(tensorLoad_1_io_tensor_rd_data_bits_0_13),
    .io_tensor_rd_data_bits_0_14(tensorLoad_1_io_tensor_rd_data_bits_0_14),
    .io_tensor_rd_data_bits_0_15(tensorLoad_1_io_tensor_rd_data_bits_0_15),
    .io_tensor_rd_data_bits_1_0(tensorLoad_1_io_tensor_rd_data_bits_1_0),
    .io_tensor_rd_data_bits_1_1(tensorLoad_1_io_tensor_rd_data_bits_1_1),
    .io_tensor_rd_data_bits_1_2(tensorLoad_1_io_tensor_rd_data_bits_1_2),
    .io_tensor_rd_data_bits_1_3(tensorLoad_1_io_tensor_rd_data_bits_1_3),
    .io_tensor_rd_data_bits_1_4(tensorLoad_1_io_tensor_rd_data_bits_1_4),
    .io_tensor_rd_data_bits_1_5(tensorLoad_1_io_tensor_rd_data_bits_1_5),
    .io_tensor_rd_data_bits_1_6(tensorLoad_1_io_tensor_rd_data_bits_1_6),
    .io_tensor_rd_data_bits_1_7(tensorLoad_1_io_tensor_rd_data_bits_1_7),
    .io_tensor_rd_data_bits_1_8(tensorLoad_1_io_tensor_rd_data_bits_1_8),
    .io_tensor_rd_data_bits_1_9(tensorLoad_1_io_tensor_rd_data_bits_1_9),
    .io_tensor_rd_data_bits_1_10(tensorLoad_1_io_tensor_rd_data_bits_1_10),
    .io_tensor_rd_data_bits_1_11(tensorLoad_1_io_tensor_rd_data_bits_1_11),
    .io_tensor_rd_data_bits_1_12(tensorLoad_1_io_tensor_rd_data_bits_1_12),
    .io_tensor_rd_data_bits_1_13(tensorLoad_1_io_tensor_rd_data_bits_1_13),
    .io_tensor_rd_data_bits_1_14(tensorLoad_1_io_tensor_rd_data_bits_1_14),
    .io_tensor_rd_data_bits_1_15(tensorLoad_1_io_tensor_rd_data_bits_1_15),
    .io_tensor_rd_data_bits_2_0(tensorLoad_1_io_tensor_rd_data_bits_2_0),
    .io_tensor_rd_data_bits_2_1(tensorLoad_1_io_tensor_rd_data_bits_2_1),
    .io_tensor_rd_data_bits_2_2(tensorLoad_1_io_tensor_rd_data_bits_2_2),
    .io_tensor_rd_data_bits_2_3(tensorLoad_1_io_tensor_rd_data_bits_2_3),
    .io_tensor_rd_data_bits_2_4(tensorLoad_1_io_tensor_rd_data_bits_2_4),
    .io_tensor_rd_data_bits_2_5(tensorLoad_1_io_tensor_rd_data_bits_2_5),
    .io_tensor_rd_data_bits_2_6(tensorLoad_1_io_tensor_rd_data_bits_2_6),
    .io_tensor_rd_data_bits_2_7(tensorLoad_1_io_tensor_rd_data_bits_2_7),
    .io_tensor_rd_data_bits_2_8(tensorLoad_1_io_tensor_rd_data_bits_2_8),
    .io_tensor_rd_data_bits_2_9(tensorLoad_1_io_tensor_rd_data_bits_2_9),
    .io_tensor_rd_data_bits_2_10(tensorLoad_1_io_tensor_rd_data_bits_2_10),
    .io_tensor_rd_data_bits_2_11(tensorLoad_1_io_tensor_rd_data_bits_2_11),
    .io_tensor_rd_data_bits_2_12(tensorLoad_1_io_tensor_rd_data_bits_2_12),
    .io_tensor_rd_data_bits_2_13(tensorLoad_1_io_tensor_rd_data_bits_2_13),
    .io_tensor_rd_data_bits_2_14(tensorLoad_1_io_tensor_rd_data_bits_2_14),
    .io_tensor_rd_data_bits_2_15(tensorLoad_1_io_tensor_rd_data_bits_2_15),
    .io_tensor_rd_data_bits_3_0(tensorLoad_1_io_tensor_rd_data_bits_3_0),
    .io_tensor_rd_data_bits_3_1(tensorLoad_1_io_tensor_rd_data_bits_3_1),
    .io_tensor_rd_data_bits_3_2(tensorLoad_1_io_tensor_rd_data_bits_3_2),
    .io_tensor_rd_data_bits_3_3(tensorLoad_1_io_tensor_rd_data_bits_3_3),
    .io_tensor_rd_data_bits_3_4(tensorLoad_1_io_tensor_rd_data_bits_3_4),
    .io_tensor_rd_data_bits_3_5(tensorLoad_1_io_tensor_rd_data_bits_3_5),
    .io_tensor_rd_data_bits_3_6(tensorLoad_1_io_tensor_rd_data_bits_3_6),
    .io_tensor_rd_data_bits_3_7(tensorLoad_1_io_tensor_rd_data_bits_3_7),
    .io_tensor_rd_data_bits_3_8(tensorLoad_1_io_tensor_rd_data_bits_3_8),
    .io_tensor_rd_data_bits_3_9(tensorLoad_1_io_tensor_rd_data_bits_3_9),
    .io_tensor_rd_data_bits_3_10(tensorLoad_1_io_tensor_rd_data_bits_3_10),
    .io_tensor_rd_data_bits_3_11(tensorLoad_1_io_tensor_rd_data_bits_3_11),
    .io_tensor_rd_data_bits_3_12(tensorLoad_1_io_tensor_rd_data_bits_3_12),
    .io_tensor_rd_data_bits_3_13(tensorLoad_1_io_tensor_rd_data_bits_3_13),
    .io_tensor_rd_data_bits_3_14(tensorLoad_1_io_tensor_rd_data_bits_3_14),
    .io_tensor_rd_data_bits_3_15(tensorLoad_1_io_tensor_rd_data_bits_3_15),
    .io_tensor_rd_data_bits_4_0(tensorLoad_1_io_tensor_rd_data_bits_4_0),
    .io_tensor_rd_data_bits_4_1(tensorLoad_1_io_tensor_rd_data_bits_4_1),
    .io_tensor_rd_data_bits_4_2(tensorLoad_1_io_tensor_rd_data_bits_4_2),
    .io_tensor_rd_data_bits_4_3(tensorLoad_1_io_tensor_rd_data_bits_4_3),
    .io_tensor_rd_data_bits_4_4(tensorLoad_1_io_tensor_rd_data_bits_4_4),
    .io_tensor_rd_data_bits_4_5(tensorLoad_1_io_tensor_rd_data_bits_4_5),
    .io_tensor_rd_data_bits_4_6(tensorLoad_1_io_tensor_rd_data_bits_4_6),
    .io_tensor_rd_data_bits_4_7(tensorLoad_1_io_tensor_rd_data_bits_4_7),
    .io_tensor_rd_data_bits_4_8(tensorLoad_1_io_tensor_rd_data_bits_4_8),
    .io_tensor_rd_data_bits_4_9(tensorLoad_1_io_tensor_rd_data_bits_4_9),
    .io_tensor_rd_data_bits_4_10(tensorLoad_1_io_tensor_rd_data_bits_4_10),
    .io_tensor_rd_data_bits_4_11(tensorLoad_1_io_tensor_rd_data_bits_4_11),
    .io_tensor_rd_data_bits_4_12(tensorLoad_1_io_tensor_rd_data_bits_4_12),
    .io_tensor_rd_data_bits_4_13(tensorLoad_1_io_tensor_rd_data_bits_4_13),
    .io_tensor_rd_data_bits_4_14(tensorLoad_1_io_tensor_rd_data_bits_4_14),
    .io_tensor_rd_data_bits_4_15(tensorLoad_1_io_tensor_rd_data_bits_4_15),
    .io_tensor_rd_data_bits_5_0(tensorLoad_1_io_tensor_rd_data_bits_5_0),
    .io_tensor_rd_data_bits_5_1(tensorLoad_1_io_tensor_rd_data_bits_5_1),
    .io_tensor_rd_data_bits_5_2(tensorLoad_1_io_tensor_rd_data_bits_5_2),
    .io_tensor_rd_data_bits_5_3(tensorLoad_1_io_tensor_rd_data_bits_5_3),
    .io_tensor_rd_data_bits_5_4(tensorLoad_1_io_tensor_rd_data_bits_5_4),
    .io_tensor_rd_data_bits_5_5(tensorLoad_1_io_tensor_rd_data_bits_5_5),
    .io_tensor_rd_data_bits_5_6(tensorLoad_1_io_tensor_rd_data_bits_5_6),
    .io_tensor_rd_data_bits_5_7(tensorLoad_1_io_tensor_rd_data_bits_5_7),
    .io_tensor_rd_data_bits_5_8(tensorLoad_1_io_tensor_rd_data_bits_5_8),
    .io_tensor_rd_data_bits_5_9(tensorLoad_1_io_tensor_rd_data_bits_5_9),
    .io_tensor_rd_data_bits_5_10(tensorLoad_1_io_tensor_rd_data_bits_5_10),
    .io_tensor_rd_data_bits_5_11(tensorLoad_1_io_tensor_rd_data_bits_5_11),
    .io_tensor_rd_data_bits_5_12(tensorLoad_1_io_tensor_rd_data_bits_5_12),
    .io_tensor_rd_data_bits_5_13(tensorLoad_1_io_tensor_rd_data_bits_5_13),
    .io_tensor_rd_data_bits_5_14(tensorLoad_1_io_tensor_rd_data_bits_5_14),
    .io_tensor_rd_data_bits_5_15(tensorLoad_1_io_tensor_rd_data_bits_5_15),
    .io_tensor_rd_data_bits_6_0(tensorLoad_1_io_tensor_rd_data_bits_6_0),
    .io_tensor_rd_data_bits_6_1(tensorLoad_1_io_tensor_rd_data_bits_6_1),
    .io_tensor_rd_data_bits_6_2(tensorLoad_1_io_tensor_rd_data_bits_6_2),
    .io_tensor_rd_data_bits_6_3(tensorLoad_1_io_tensor_rd_data_bits_6_3),
    .io_tensor_rd_data_bits_6_4(tensorLoad_1_io_tensor_rd_data_bits_6_4),
    .io_tensor_rd_data_bits_6_5(tensorLoad_1_io_tensor_rd_data_bits_6_5),
    .io_tensor_rd_data_bits_6_6(tensorLoad_1_io_tensor_rd_data_bits_6_6),
    .io_tensor_rd_data_bits_6_7(tensorLoad_1_io_tensor_rd_data_bits_6_7),
    .io_tensor_rd_data_bits_6_8(tensorLoad_1_io_tensor_rd_data_bits_6_8),
    .io_tensor_rd_data_bits_6_9(tensorLoad_1_io_tensor_rd_data_bits_6_9),
    .io_tensor_rd_data_bits_6_10(tensorLoad_1_io_tensor_rd_data_bits_6_10),
    .io_tensor_rd_data_bits_6_11(tensorLoad_1_io_tensor_rd_data_bits_6_11),
    .io_tensor_rd_data_bits_6_12(tensorLoad_1_io_tensor_rd_data_bits_6_12),
    .io_tensor_rd_data_bits_6_13(tensorLoad_1_io_tensor_rd_data_bits_6_13),
    .io_tensor_rd_data_bits_6_14(tensorLoad_1_io_tensor_rd_data_bits_6_14),
    .io_tensor_rd_data_bits_6_15(tensorLoad_1_io_tensor_rd_data_bits_6_15),
    .io_tensor_rd_data_bits_7_0(tensorLoad_1_io_tensor_rd_data_bits_7_0),
    .io_tensor_rd_data_bits_7_1(tensorLoad_1_io_tensor_rd_data_bits_7_1),
    .io_tensor_rd_data_bits_7_2(tensorLoad_1_io_tensor_rd_data_bits_7_2),
    .io_tensor_rd_data_bits_7_3(tensorLoad_1_io_tensor_rd_data_bits_7_3),
    .io_tensor_rd_data_bits_7_4(tensorLoad_1_io_tensor_rd_data_bits_7_4),
    .io_tensor_rd_data_bits_7_5(tensorLoad_1_io_tensor_rd_data_bits_7_5),
    .io_tensor_rd_data_bits_7_6(tensorLoad_1_io_tensor_rd_data_bits_7_6),
    .io_tensor_rd_data_bits_7_7(tensorLoad_1_io_tensor_rd_data_bits_7_7),
    .io_tensor_rd_data_bits_7_8(tensorLoad_1_io_tensor_rd_data_bits_7_8),
    .io_tensor_rd_data_bits_7_9(tensorLoad_1_io_tensor_rd_data_bits_7_9),
    .io_tensor_rd_data_bits_7_10(tensorLoad_1_io_tensor_rd_data_bits_7_10),
    .io_tensor_rd_data_bits_7_11(tensorLoad_1_io_tensor_rd_data_bits_7_11),
    .io_tensor_rd_data_bits_7_12(tensorLoad_1_io_tensor_rd_data_bits_7_12),
    .io_tensor_rd_data_bits_7_13(tensorLoad_1_io_tensor_rd_data_bits_7_13),
    .io_tensor_rd_data_bits_7_14(tensorLoad_1_io_tensor_rd_data_bits_7_14),
    .io_tensor_rd_data_bits_7_15(tensorLoad_1_io_tensor_rd_data_bits_7_15),
    .io_tensor_rd_data_bits_8_0(tensorLoad_1_io_tensor_rd_data_bits_8_0),
    .io_tensor_rd_data_bits_8_1(tensorLoad_1_io_tensor_rd_data_bits_8_1),
    .io_tensor_rd_data_bits_8_2(tensorLoad_1_io_tensor_rd_data_bits_8_2),
    .io_tensor_rd_data_bits_8_3(tensorLoad_1_io_tensor_rd_data_bits_8_3),
    .io_tensor_rd_data_bits_8_4(tensorLoad_1_io_tensor_rd_data_bits_8_4),
    .io_tensor_rd_data_bits_8_5(tensorLoad_1_io_tensor_rd_data_bits_8_5),
    .io_tensor_rd_data_bits_8_6(tensorLoad_1_io_tensor_rd_data_bits_8_6),
    .io_tensor_rd_data_bits_8_7(tensorLoad_1_io_tensor_rd_data_bits_8_7),
    .io_tensor_rd_data_bits_8_8(tensorLoad_1_io_tensor_rd_data_bits_8_8),
    .io_tensor_rd_data_bits_8_9(tensorLoad_1_io_tensor_rd_data_bits_8_9),
    .io_tensor_rd_data_bits_8_10(tensorLoad_1_io_tensor_rd_data_bits_8_10),
    .io_tensor_rd_data_bits_8_11(tensorLoad_1_io_tensor_rd_data_bits_8_11),
    .io_tensor_rd_data_bits_8_12(tensorLoad_1_io_tensor_rd_data_bits_8_12),
    .io_tensor_rd_data_bits_8_13(tensorLoad_1_io_tensor_rd_data_bits_8_13),
    .io_tensor_rd_data_bits_8_14(tensorLoad_1_io_tensor_rd_data_bits_8_14),
    .io_tensor_rd_data_bits_8_15(tensorLoad_1_io_tensor_rd_data_bits_8_15),
    .io_tensor_rd_data_bits_9_0(tensorLoad_1_io_tensor_rd_data_bits_9_0),
    .io_tensor_rd_data_bits_9_1(tensorLoad_1_io_tensor_rd_data_bits_9_1),
    .io_tensor_rd_data_bits_9_2(tensorLoad_1_io_tensor_rd_data_bits_9_2),
    .io_tensor_rd_data_bits_9_3(tensorLoad_1_io_tensor_rd_data_bits_9_3),
    .io_tensor_rd_data_bits_9_4(tensorLoad_1_io_tensor_rd_data_bits_9_4),
    .io_tensor_rd_data_bits_9_5(tensorLoad_1_io_tensor_rd_data_bits_9_5),
    .io_tensor_rd_data_bits_9_6(tensorLoad_1_io_tensor_rd_data_bits_9_6),
    .io_tensor_rd_data_bits_9_7(tensorLoad_1_io_tensor_rd_data_bits_9_7),
    .io_tensor_rd_data_bits_9_8(tensorLoad_1_io_tensor_rd_data_bits_9_8),
    .io_tensor_rd_data_bits_9_9(tensorLoad_1_io_tensor_rd_data_bits_9_9),
    .io_tensor_rd_data_bits_9_10(tensorLoad_1_io_tensor_rd_data_bits_9_10),
    .io_tensor_rd_data_bits_9_11(tensorLoad_1_io_tensor_rd_data_bits_9_11),
    .io_tensor_rd_data_bits_9_12(tensorLoad_1_io_tensor_rd_data_bits_9_12),
    .io_tensor_rd_data_bits_9_13(tensorLoad_1_io_tensor_rd_data_bits_9_13),
    .io_tensor_rd_data_bits_9_14(tensorLoad_1_io_tensor_rd_data_bits_9_14),
    .io_tensor_rd_data_bits_9_15(tensorLoad_1_io_tensor_rd_data_bits_9_15),
    .io_tensor_rd_data_bits_10_0(tensorLoad_1_io_tensor_rd_data_bits_10_0),
    .io_tensor_rd_data_bits_10_1(tensorLoad_1_io_tensor_rd_data_bits_10_1),
    .io_tensor_rd_data_bits_10_2(tensorLoad_1_io_tensor_rd_data_bits_10_2),
    .io_tensor_rd_data_bits_10_3(tensorLoad_1_io_tensor_rd_data_bits_10_3),
    .io_tensor_rd_data_bits_10_4(tensorLoad_1_io_tensor_rd_data_bits_10_4),
    .io_tensor_rd_data_bits_10_5(tensorLoad_1_io_tensor_rd_data_bits_10_5),
    .io_tensor_rd_data_bits_10_6(tensorLoad_1_io_tensor_rd_data_bits_10_6),
    .io_tensor_rd_data_bits_10_7(tensorLoad_1_io_tensor_rd_data_bits_10_7),
    .io_tensor_rd_data_bits_10_8(tensorLoad_1_io_tensor_rd_data_bits_10_8),
    .io_tensor_rd_data_bits_10_9(tensorLoad_1_io_tensor_rd_data_bits_10_9),
    .io_tensor_rd_data_bits_10_10(tensorLoad_1_io_tensor_rd_data_bits_10_10),
    .io_tensor_rd_data_bits_10_11(tensorLoad_1_io_tensor_rd_data_bits_10_11),
    .io_tensor_rd_data_bits_10_12(tensorLoad_1_io_tensor_rd_data_bits_10_12),
    .io_tensor_rd_data_bits_10_13(tensorLoad_1_io_tensor_rd_data_bits_10_13),
    .io_tensor_rd_data_bits_10_14(tensorLoad_1_io_tensor_rd_data_bits_10_14),
    .io_tensor_rd_data_bits_10_15(tensorLoad_1_io_tensor_rd_data_bits_10_15),
    .io_tensor_rd_data_bits_11_0(tensorLoad_1_io_tensor_rd_data_bits_11_0),
    .io_tensor_rd_data_bits_11_1(tensorLoad_1_io_tensor_rd_data_bits_11_1),
    .io_tensor_rd_data_bits_11_2(tensorLoad_1_io_tensor_rd_data_bits_11_2),
    .io_tensor_rd_data_bits_11_3(tensorLoad_1_io_tensor_rd_data_bits_11_3),
    .io_tensor_rd_data_bits_11_4(tensorLoad_1_io_tensor_rd_data_bits_11_4),
    .io_tensor_rd_data_bits_11_5(tensorLoad_1_io_tensor_rd_data_bits_11_5),
    .io_tensor_rd_data_bits_11_6(tensorLoad_1_io_tensor_rd_data_bits_11_6),
    .io_tensor_rd_data_bits_11_7(tensorLoad_1_io_tensor_rd_data_bits_11_7),
    .io_tensor_rd_data_bits_11_8(tensorLoad_1_io_tensor_rd_data_bits_11_8),
    .io_tensor_rd_data_bits_11_9(tensorLoad_1_io_tensor_rd_data_bits_11_9),
    .io_tensor_rd_data_bits_11_10(tensorLoad_1_io_tensor_rd_data_bits_11_10),
    .io_tensor_rd_data_bits_11_11(tensorLoad_1_io_tensor_rd_data_bits_11_11),
    .io_tensor_rd_data_bits_11_12(tensorLoad_1_io_tensor_rd_data_bits_11_12),
    .io_tensor_rd_data_bits_11_13(tensorLoad_1_io_tensor_rd_data_bits_11_13),
    .io_tensor_rd_data_bits_11_14(tensorLoad_1_io_tensor_rd_data_bits_11_14),
    .io_tensor_rd_data_bits_11_15(tensorLoad_1_io_tensor_rd_data_bits_11_15),
    .io_tensor_rd_data_bits_12_0(tensorLoad_1_io_tensor_rd_data_bits_12_0),
    .io_tensor_rd_data_bits_12_1(tensorLoad_1_io_tensor_rd_data_bits_12_1),
    .io_tensor_rd_data_bits_12_2(tensorLoad_1_io_tensor_rd_data_bits_12_2),
    .io_tensor_rd_data_bits_12_3(tensorLoad_1_io_tensor_rd_data_bits_12_3),
    .io_tensor_rd_data_bits_12_4(tensorLoad_1_io_tensor_rd_data_bits_12_4),
    .io_tensor_rd_data_bits_12_5(tensorLoad_1_io_tensor_rd_data_bits_12_5),
    .io_tensor_rd_data_bits_12_6(tensorLoad_1_io_tensor_rd_data_bits_12_6),
    .io_tensor_rd_data_bits_12_7(tensorLoad_1_io_tensor_rd_data_bits_12_7),
    .io_tensor_rd_data_bits_12_8(tensorLoad_1_io_tensor_rd_data_bits_12_8),
    .io_tensor_rd_data_bits_12_9(tensorLoad_1_io_tensor_rd_data_bits_12_9),
    .io_tensor_rd_data_bits_12_10(tensorLoad_1_io_tensor_rd_data_bits_12_10),
    .io_tensor_rd_data_bits_12_11(tensorLoad_1_io_tensor_rd_data_bits_12_11),
    .io_tensor_rd_data_bits_12_12(tensorLoad_1_io_tensor_rd_data_bits_12_12),
    .io_tensor_rd_data_bits_12_13(tensorLoad_1_io_tensor_rd_data_bits_12_13),
    .io_tensor_rd_data_bits_12_14(tensorLoad_1_io_tensor_rd_data_bits_12_14),
    .io_tensor_rd_data_bits_12_15(tensorLoad_1_io_tensor_rd_data_bits_12_15),
    .io_tensor_rd_data_bits_13_0(tensorLoad_1_io_tensor_rd_data_bits_13_0),
    .io_tensor_rd_data_bits_13_1(tensorLoad_1_io_tensor_rd_data_bits_13_1),
    .io_tensor_rd_data_bits_13_2(tensorLoad_1_io_tensor_rd_data_bits_13_2),
    .io_tensor_rd_data_bits_13_3(tensorLoad_1_io_tensor_rd_data_bits_13_3),
    .io_tensor_rd_data_bits_13_4(tensorLoad_1_io_tensor_rd_data_bits_13_4),
    .io_tensor_rd_data_bits_13_5(tensorLoad_1_io_tensor_rd_data_bits_13_5),
    .io_tensor_rd_data_bits_13_6(tensorLoad_1_io_tensor_rd_data_bits_13_6),
    .io_tensor_rd_data_bits_13_7(tensorLoad_1_io_tensor_rd_data_bits_13_7),
    .io_tensor_rd_data_bits_13_8(tensorLoad_1_io_tensor_rd_data_bits_13_8),
    .io_tensor_rd_data_bits_13_9(tensorLoad_1_io_tensor_rd_data_bits_13_9),
    .io_tensor_rd_data_bits_13_10(tensorLoad_1_io_tensor_rd_data_bits_13_10),
    .io_tensor_rd_data_bits_13_11(tensorLoad_1_io_tensor_rd_data_bits_13_11),
    .io_tensor_rd_data_bits_13_12(tensorLoad_1_io_tensor_rd_data_bits_13_12),
    .io_tensor_rd_data_bits_13_13(tensorLoad_1_io_tensor_rd_data_bits_13_13),
    .io_tensor_rd_data_bits_13_14(tensorLoad_1_io_tensor_rd_data_bits_13_14),
    .io_tensor_rd_data_bits_13_15(tensorLoad_1_io_tensor_rd_data_bits_13_15),
    .io_tensor_rd_data_bits_14_0(tensorLoad_1_io_tensor_rd_data_bits_14_0),
    .io_tensor_rd_data_bits_14_1(tensorLoad_1_io_tensor_rd_data_bits_14_1),
    .io_tensor_rd_data_bits_14_2(tensorLoad_1_io_tensor_rd_data_bits_14_2),
    .io_tensor_rd_data_bits_14_3(tensorLoad_1_io_tensor_rd_data_bits_14_3),
    .io_tensor_rd_data_bits_14_4(tensorLoad_1_io_tensor_rd_data_bits_14_4),
    .io_tensor_rd_data_bits_14_5(tensorLoad_1_io_tensor_rd_data_bits_14_5),
    .io_tensor_rd_data_bits_14_6(tensorLoad_1_io_tensor_rd_data_bits_14_6),
    .io_tensor_rd_data_bits_14_7(tensorLoad_1_io_tensor_rd_data_bits_14_7),
    .io_tensor_rd_data_bits_14_8(tensorLoad_1_io_tensor_rd_data_bits_14_8),
    .io_tensor_rd_data_bits_14_9(tensorLoad_1_io_tensor_rd_data_bits_14_9),
    .io_tensor_rd_data_bits_14_10(tensorLoad_1_io_tensor_rd_data_bits_14_10),
    .io_tensor_rd_data_bits_14_11(tensorLoad_1_io_tensor_rd_data_bits_14_11),
    .io_tensor_rd_data_bits_14_12(tensorLoad_1_io_tensor_rd_data_bits_14_12),
    .io_tensor_rd_data_bits_14_13(tensorLoad_1_io_tensor_rd_data_bits_14_13),
    .io_tensor_rd_data_bits_14_14(tensorLoad_1_io_tensor_rd_data_bits_14_14),
    .io_tensor_rd_data_bits_14_15(tensorLoad_1_io_tensor_rd_data_bits_14_15),
    .io_tensor_rd_data_bits_15_0(tensorLoad_1_io_tensor_rd_data_bits_15_0),
    .io_tensor_rd_data_bits_15_1(tensorLoad_1_io_tensor_rd_data_bits_15_1),
    .io_tensor_rd_data_bits_15_2(tensorLoad_1_io_tensor_rd_data_bits_15_2),
    .io_tensor_rd_data_bits_15_3(tensorLoad_1_io_tensor_rd_data_bits_15_3),
    .io_tensor_rd_data_bits_15_4(tensorLoad_1_io_tensor_rd_data_bits_15_4),
    .io_tensor_rd_data_bits_15_5(tensorLoad_1_io_tensor_rd_data_bits_15_5),
    .io_tensor_rd_data_bits_15_6(tensorLoad_1_io_tensor_rd_data_bits_15_6),
    .io_tensor_rd_data_bits_15_7(tensorLoad_1_io_tensor_rd_data_bits_15_7),
    .io_tensor_rd_data_bits_15_8(tensorLoad_1_io_tensor_rd_data_bits_15_8),
    .io_tensor_rd_data_bits_15_9(tensorLoad_1_io_tensor_rd_data_bits_15_9),
    .io_tensor_rd_data_bits_15_10(tensorLoad_1_io_tensor_rd_data_bits_15_10),
    .io_tensor_rd_data_bits_15_11(tensorLoad_1_io_tensor_rd_data_bits_15_11),
    .io_tensor_rd_data_bits_15_12(tensorLoad_1_io_tensor_rd_data_bits_15_12),
    .io_tensor_rd_data_bits_15_13(tensorLoad_1_io_tensor_rd_data_bits_15_13),
    .io_tensor_rd_data_bits_15_14(tensorLoad_1_io_tensor_rd_data_bits_15_14),
    .io_tensor_rd_data_bits_15_15(tensorLoad_1_io_tensor_rd_data_bits_15_15)
  );
  assign _T_4999 = dec_io_pop_next ? s_io_sready : 1'h1; // @[Load.scala 60:40:@5320.4]
  assign start = inst_q_io_deq_valid & _T_4999; // @[Load.scala 60:35:@5321.4]
  assign done = dec_io_isInput ? tensorLoad_0_io_done : tensorLoad_1_io_done; // @[Load.scala 61:17:@5322.4]
  assign _T_5000 = 2'h0 == state; // @[Conditional.scala 37:30:@5323.4]
  assign _T_5001 = dec_io_isInput | dec_io_isWeight; // @[Load.scala 69:35:@5330.10]
  assign _GEN_0 = _T_5001 ? 2'h2 : state; // @[Load.scala 69:55:@5331.10]
  assign _GEN_1 = dec_io_isSync ? 2'h1 : _GEN_0; // @[Load.scala 67:29:@5326.8]
  assign _GEN_2 = start ? _GEN_1 : state; // @[Load.scala 66:19:@5325.6]
  assign _T_5002 = 2'h1 == state; // @[Conditional.scala 37:30:@5337.6]
  assign _T_5003 = 2'h2 == state; // @[Conditional.scala 37:30:@5342.8]
  assign _GEN_3 = done ? 2'h0 : state; // @[Load.scala 78:18:@5344.10]
  assign _GEN_4 = _T_5003 ? _GEN_3 : state; // @[Conditional.scala 39:67:@5343.8]
  assign _GEN_5 = _T_5002 ? 2'h0 : _GEN_4; // @[Conditional.scala 39:67:@5338.6]
  assign _GEN_6 = _T_5000 ? _GEN_2 : _GEN_5; // @[Conditional.scala 40:58:@5324.4]
  assign _T_5004 = state == 2'h2; // @[Load.scala 86:33:@5351.4]
  assign _T_5005 = _T_5004 & done; // @[Load.scala 86:42:@5352.4]
  assign _T_5006 = state == 2'h1; // @[Load.scala 86:59:@5353.4]
  assign _T_5007 = _T_5005 | _T_5006; // @[Load.scala 86:50:@5354.4]
  assign _T_5008 = state == 2'h0; // @[Load.scala 94:37:@5356.4]
  assign _T_5009 = _T_5008 & start; // @[Load.scala 94:47:@5357.4]
  assign io_o_post = dec_io_push_next & _T_5007; // @[Load.scala 104:13:@5946.4]
  assign io_inst_ready = inst_q_io_enq_ready; // @[Load.scala 85:17:@5350.4]
  assign io_vme_rd_0_cmd_valid = tensorLoad_0_io_vme_rd_cmd_valid; // @[Load.scala 98:18:@5404.4]
  assign io_vme_rd_0_cmd_bits_addr = tensorLoad_0_io_vme_rd_cmd_bits_addr; // @[Load.scala 98:18:@5403.4]
  assign io_vme_rd_0_cmd_bits_len = tensorLoad_0_io_vme_rd_cmd_bits_len; // @[Load.scala 98:18:@5402.4]
  assign io_vme_rd_0_data_ready = tensorLoad_0_io_vme_rd_data_ready; // @[Load.scala 98:18:@5401.4]
  assign io_vme_rd_1_cmd_valid = tensorLoad_1_io_vme_rd_cmd_valid; // @[Load.scala 98:18:@5934.4]
  assign io_vme_rd_1_cmd_bits_addr = tensorLoad_1_io_vme_rd_cmd_bits_addr; // @[Load.scala 98:18:@5933.4]
  assign io_vme_rd_1_cmd_bits_len = tensorLoad_1_io_vme_rd_cmd_bits_len; // @[Load.scala 98:18:@5932.4]
  assign io_vme_rd_1_data_ready = tensorLoad_1_io_vme_rd_data_ready; // @[Load.scala 98:18:@5931.4]
  assign io_inp_rd_data_valid = tensorLoad_0_io_tensor_rd_data_valid; // @[Load.scala 97:29:@5396.4]
  assign io_inp_rd_data_bits_0_0 = tensorLoad_0_io_tensor_rd_data_bits_0_0; // @[Load.scala 97:29:@5380.4]
  assign io_inp_rd_data_bits_0_1 = tensorLoad_0_io_tensor_rd_data_bits_0_1; // @[Load.scala 97:29:@5381.4]
  assign io_inp_rd_data_bits_0_2 = tensorLoad_0_io_tensor_rd_data_bits_0_2; // @[Load.scala 97:29:@5382.4]
  assign io_inp_rd_data_bits_0_3 = tensorLoad_0_io_tensor_rd_data_bits_0_3; // @[Load.scala 97:29:@5383.4]
  assign io_inp_rd_data_bits_0_4 = tensorLoad_0_io_tensor_rd_data_bits_0_4; // @[Load.scala 97:29:@5384.4]
  assign io_inp_rd_data_bits_0_5 = tensorLoad_0_io_tensor_rd_data_bits_0_5; // @[Load.scala 97:29:@5385.4]
  assign io_inp_rd_data_bits_0_6 = tensorLoad_0_io_tensor_rd_data_bits_0_6; // @[Load.scala 97:29:@5386.4]
  assign io_inp_rd_data_bits_0_7 = tensorLoad_0_io_tensor_rd_data_bits_0_7; // @[Load.scala 97:29:@5387.4]
  assign io_inp_rd_data_bits_0_8 = tensorLoad_0_io_tensor_rd_data_bits_0_8; // @[Load.scala 97:29:@5388.4]
  assign io_inp_rd_data_bits_0_9 = tensorLoad_0_io_tensor_rd_data_bits_0_9; // @[Load.scala 97:29:@5389.4]
  assign io_inp_rd_data_bits_0_10 = tensorLoad_0_io_tensor_rd_data_bits_0_10; // @[Load.scala 97:29:@5390.4]
  assign io_inp_rd_data_bits_0_11 = tensorLoad_0_io_tensor_rd_data_bits_0_11; // @[Load.scala 97:29:@5391.4]
  assign io_inp_rd_data_bits_0_12 = tensorLoad_0_io_tensor_rd_data_bits_0_12; // @[Load.scala 97:29:@5392.4]
  assign io_inp_rd_data_bits_0_13 = tensorLoad_0_io_tensor_rd_data_bits_0_13; // @[Load.scala 97:29:@5393.4]
  assign io_inp_rd_data_bits_0_14 = tensorLoad_0_io_tensor_rd_data_bits_0_14; // @[Load.scala 97:29:@5394.4]
  assign io_inp_rd_data_bits_0_15 = tensorLoad_0_io_tensor_rd_data_bits_0_15; // @[Load.scala 97:29:@5395.4]
  assign io_wgt_rd_data_valid = tensorLoad_1_io_tensor_rd_data_valid; // @[Load.scala 97:29:@5926.4]
  assign io_wgt_rd_data_bits_0_0 = tensorLoad_1_io_tensor_rd_data_bits_0_0; // @[Load.scala 97:29:@5670.4]
  assign io_wgt_rd_data_bits_0_1 = tensorLoad_1_io_tensor_rd_data_bits_0_1; // @[Load.scala 97:29:@5671.4]
  assign io_wgt_rd_data_bits_0_2 = tensorLoad_1_io_tensor_rd_data_bits_0_2; // @[Load.scala 97:29:@5672.4]
  assign io_wgt_rd_data_bits_0_3 = tensorLoad_1_io_tensor_rd_data_bits_0_3; // @[Load.scala 97:29:@5673.4]
  assign io_wgt_rd_data_bits_0_4 = tensorLoad_1_io_tensor_rd_data_bits_0_4; // @[Load.scala 97:29:@5674.4]
  assign io_wgt_rd_data_bits_0_5 = tensorLoad_1_io_tensor_rd_data_bits_0_5; // @[Load.scala 97:29:@5675.4]
  assign io_wgt_rd_data_bits_0_6 = tensorLoad_1_io_tensor_rd_data_bits_0_6; // @[Load.scala 97:29:@5676.4]
  assign io_wgt_rd_data_bits_0_7 = tensorLoad_1_io_tensor_rd_data_bits_0_7; // @[Load.scala 97:29:@5677.4]
  assign io_wgt_rd_data_bits_0_8 = tensorLoad_1_io_tensor_rd_data_bits_0_8; // @[Load.scala 97:29:@5678.4]
  assign io_wgt_rd_data_bits_0_9 = tensorLoad_1_io_tensor_rd_data_bits_0_9; // @[Load.scala 97:29:@5679.4]
  assign io_wgt_rd_data_bits_0_10 = tensorLoad_1_io_tensor_rd_data_bits_0_10; // @[Load.scala 97:29:@5680.4]
  assign io_wgt_rd_data_bits_0_11 = tensorLoad_1_io_tensor_rd_data_bits_0_11; // @[Load.scala 97:29:@5681.4]
  assign io_wgt_rd_data_bits_0_12 = tensorLoad_1_io_tensor_rd_data_bits_0_12; // @[Load.scala 97:29:@5682.4]
  assign io_wgt_rd_data_bits_0_13 = tensorLoad_1_io_tensor_rd_data_bits_0_13; // @[Load.scala 97:29:@5683.4]
  assign io_wgt_rd_data_bits_0_14 = tensorLoad_1_io_tensor_rd_data_bits_0_14; // @[Load.scala 97:29:@5684.4]
  assign io_wgt_rd_data_bits_0_15 = tensorLoad_1_io_tensor_rd_data_bits_0_15; // @[Load.scala 97:29:@5685.4]
  assign io_wgt_rd_data_bits_1_0 = tensorLoad_1_io_tensor_rd_data_bits_1_0; // @[Load.scala 97:29:@5686.4]
  assign io_wgt_rd_data_bits_1_1 = tensorLoad_1_io_tensor_rd_data_bits_1_1; // @[Load.scala 97:29:@5687.4]
  assign io_wgt_rd_data_bits_1_2 = tensorLoad_1_io_tensor_rd_data_bits_1_2; // @[Load.scala 97:29:@5688.4]
  assign io_wgt_rd_data_bits_1_3 = tensorLoad_1_io_tensor_rd_data_bits_1_3; // @[Load.scala 97:29:@5689.4]
  assign io_wgt_rd_data_bits_1_4 = tensorLoad_1_io_tensor_rd_data_bits_1_4; // @[Load.scala 97:29:@5690.4]
  assign io_wgt_rd_data_bits_1_5 = tensorLoad_1_io_tensor_rd_data_bits_1_5; // @[Load.scala 97:29:@5691.4]
  assign io_wgt_rd_data_bits_1_6 = tensorLoad_1_io_tensor_rd_data_bits_1_6; // @[Load.scala 97:29:@5692.4]
  assign io_wgt_rd_data_bits_1_7 = tensorLoad_1_io_tensor_rd_data_bits_1_7; // @[Load.scala 97:29:@5693.4]
  assign io_wgt_rd_data_bits_1_8 = tensorLoad_1_io_tensor_rd_data_bits_1_8; // @[Load.scala 97:29:@5694.4]
  assign io_wgt_rd_data_bits_1_9 = tensorLoad_1_io_tensor_rd_data_bits_1_9; // @[Load.scala 97:29:@5695.4]
  assign io_wgt_rd_data_bits_1_10 = tensorLoad_1_io_tensor_rd_data_bits_1_10; // @[Load.scala 97:29:@5696.4]
  assign io_wgt_rd_data_bits_1_11 = tensorLoad_1_io_tensor_rd_data_bits_1_11; // @[Load.scala 97:29:@5697.4]
  assign io_wgt_rd_data_bits_1_12 = tensorLoad_1_io_tensor_rd_data_bits_1_12; // @[Load.scala 97:29:@5698.4]
  assign io_wgt_rd_data_bits_1_13 = tensorLoad_1_io_tensor_rd_data_bits_1_13; // @[Load.scala 97:29:@5699.4]
  assign io_wgt_rd_data_bits_1_14 = tensorLoad_1_io_tensor_rd_data_bits_1_14; // @[Load.scala 97:29:@5700.4]
  assign io_wgt_rd_data_bits_1_15 = tensorLoad_1_io_tensor_rd_data_bits_1_15; // @[Load.scala 97:29:@5701.4]
  assign io_wgt_rd_data_bits_2_0 = tensorLoad_1_io_tensor_rd_data_bits_2_0; // @[Load.scala 97:29:@5702.4]
  assign io_wgt_rd_data_bits_2_1 = tensorLoad_1_io_tensor_rd_data_bits_2_1; // @[Load.scala 97:29:@5703.4]
  assign io_wgt_rd_data_bits_2_2 = tensorLoad_1_io_tensor_rd_data_bits_2_2; // @[Load.scala 97:29:@5704.4]
  assign io_wgt_rd_data_bits_2_3 = tensorLoad_1_io_tensor_rd_data_bits_2_3; // @[Load.scala 97:29:@5705.4]
  assign io_wgt_rd_data_bits_2_4 = tensorLoad_1_io_tensor_rd_data_bits_2_4; // @[Load.scala 97:29:@5706.4]
  assign io_wgt_rd_data_bits_2_5 = tensorLoad_1_io_tensor_rd_data_bits_2_5; // @[Load.scala 97:29:@5707.4]
  assign io_wgt_rd_data_bits_2_6 = tensorLoad_1_io_tensor_rd_data_bits_2_6; // @[Load.scala 97:29:@5708.4]
  assign io_wgt_rd_data_bits_2_7 = tensorLoad_1_io_tensor_rd_data_bits_2_7; // @[Load.scala 97:29:@5709.4]
  assign io_wgt_rd_data_bits_2_8 = tensorLoad_1_io_tensor_rd_data_bits_2_8; // @[Load.scala 97:29:@5710.4]
  assign io_wgt_rd_data_bits_2_9 = tensorLoad_1_io_tensor_rd_data_bits_2_9; // @[Load.scala 97:29:@5711.4]
  assign io_wgt_rd_data_bits_2_10 = tensorLoad_1_io_tensor_rd_data_bits_2_10; // @[Load.scala 97:29:@5712.4]
  assign io_wgt_rd_data_bits_2_11 = tensorLoad_1_io_tensor_rd_data_bits_2_11; // @[Load.scala 97:29:@5713.4]
  assign io_wgt_rd_data_bits_2_12 = tensorLoad_1_io_tensor_rd_data_bits_2_12; // @[Load.scala 97:29:@5714.4]
  assign io_wgt_rd_data_bits_2_13 = tensorLoad_1_io_tensor_rd_data_bits_2_13; // @[Load.scala 97:29:@5715.4]
  assign io_wgt_rd_data_bits_2_14 = tensorLoad_1_io_tensor_rd_data_bits_2_14; // @[Load.scala 97:29:@5716.4]
  assign io_wgt_rd_data_bits_2_15 = tensorLoad_1_io_tensor_rd_data_bits_2_15; // @[Load.scala 97:29:@5717.4]
  assign io_wgt_rd_data_bits_3_0 = tensorLoad_1_io_tensor_rd_data_bits_3_0; // @[Load.scala 97:29:@5718.4]
  assign io_wgt_rd_data_bits_3_1 = tensorLoad_1_io_tensor_rd_data_bits_3_1; // @[Load.scala 97:29:@5719.4]
  assign io_wgt_rd_data_bits_3_2 = tensorLoad_1_io_tensor_rd_data_bits_3_2; // @[Load.scala 97:29:@5720.4]
  assign io_wgt_rd_data_bits_3_3 = tensorLoad_1_io_tensor_rd_data_bits_3_3; // @[Load.scala 97:29:@5721.4]
  assign io_wgt_rd_data_bits_3_4 = tensorLoad_1_io_tensor_rd_data_bits_3_4; // @[Load.scala 97:29:@5722.4]
  assign io_wgt_rd_data_bits_3_5 = tensorLoad_1_io_tensor_rd_data_bits_3_5; // @[Load.scala 97:29:@5723.4]
  assign io_wgt_rd_data_bits_3_6 = tensorLoad_1_io_tensor_rd_data_bits_3_6; // @[Load.scala 97:29:@5724.4]
  assign io_wgt_rd_data_bits_3_7 = tensorLoad_1_io_tensor_rd_data_bits_3_7; // @[Load.scala 97:29:@5725.4]
  assign io_wgt_rd_data_bits_3_8 = tensorLoad_1_io_tensor_rd_data_bits_3_8; // @[Load.scala 97:29:@5726.4]
  assign io_wgt_rd_data_bits_3_9 = tensorLoad_1_io_tensor_rd_data_bits_3_9; // @[Load.scala 97:29:@5727.4]
  assign io_wgt_rd_data_bits_3_10 = tensorLoad_1_io_tensor_rd_data_bits_3_10; // @[Load.scala 97:29:@5728.4]
  assign io_wgt_rd_data_bits_3_11 = tensorLoad_1_io_tensor_rd_data_bits_3_11; // @[Load.scala 97:29:@5729.4]
  assign io_wgt_rd_data_bits_3_12 = tensorLoad_1_io_tensor_rd_data_bits_3_12; // @[Load.scala 97:29:@5730.4]
  assign io_wgt_rd_data_bits_3_13 = tensorLoad_1_io_tensor_rd_data_bits_3_13; // @[Load.scala 97:29:@5731.4]
  assign io_wgt_rd_data_bits_3_14 = tensorLoad_1_io_tensor_rd_data_bits_3_14; // @[Load.scala 97:29:@5732.4]
  assign io_wgt_rd_data_bits_3_15 = tensorLoad_1_io_tensor_rd_data_bits_3_15; // @[Load.scala 97:29:@5733.4]
  assign io_wgt_rd_data_bits_4_0 = tensorLoad_1_io_tensor_rd_data_bits_4_0; // @[Load.scala 97:29:@5734.4]
  assign io_wgt_rd_data_bits_4_1 = tensorLoad_1_io_tensor_rd_data_bits_4_1; // @[Load.scala 97:29:@5735.4]
  assign io_wgt_rd_data_bits_4_2 = tensorLoad_1_io_tensor_rd_data_bits_4_2; // @[Load.scala 97:29:@5736.4]
  assign io_wgt_rd_data_bits_4_3 = tensorLoad_1_io_tensor_rd_data_bits_4_3; // @[Load.scala 97:29:@5737.4]
  assign io_wgt_rd_data_bits_4_4 = tensorLoad_1_io_tensor_rd_data_bits_4_4; // @[Load.scala 97:29:@5738.4]
  assign io_wgt_rd_data_bits_4_5 = tensorLoad_1_io_tensor_rd_data_bits_4_5; // @[Load.scala 97:29:@5739.4]
  assign io_wgt_rd_data_bits_4_6 = tensorLoad_1_io_tensor_rd_data_bits_4_6; // @[Load.scala 97:29:@5740.4]
  assign io_wgt_rd_data_bits_4_7 = tensorLoad_1_io_tensor_rd_data_bits_4_7; // @[Load.scala 97:29:@5741.4]
  assign io_wgt_rd_data_bits_4_8 = tensorLoad_1_io_tensor_rd_data_bits_4_8; // @[Load.scala 97:29:@5742.4]
  assign io_wgt_rd_data_bits_4_9 = tensorLoad_1_io_tensor_rd_data_bits_4_9; // @[Load.scala 97:29:@5743.4]
  assign io_wgt_rd_data_bits_4_10 = tensorLoad_1_io_tensor_rd_data_bits_4_10; // @[Load.scala 97:29:@5744.4]
  assign io_wgt_rd_data_bits_4_11 = tensorLoad_1_io_tensor_rd_data_bits_4_11; // @[Load.scala 97:29:@5745.4]
  assign io_wgt_rd_data_bits_4_12 = tensorLoad_1_io_tensor_rd_data_bits_4_12; // @[Load.scala 97:29:@5746.4]
  assign io_wgt_rd_data_bits_4_13 = tensorLoad_1_io_tensor_rd_data_bits_4_13; // @[Load.scala 97:29:@5747.4]
  assign io_wgt_rd_data_bits_4_14 = tensorLoad_1_io_tensor_rd_data_bits_4_14; // @[Load.scala 97:29:@5748.4]
  assign io_wgt_rd_data_bits_4_15 = tensorLoad_1_io_tensor_rd_data_bits_4_15; // @[Load.scala 97:29:@5749.4]
  assign io_wgt_rd_data_bits_5_0 = tensorLoad_1_io_tensor_rd_data_bits_5_0; // @[Load.scala 97:29:@5750.4]
  assign io_wgt_rd_data_bits_5_1 = tensorLoad_1_io_tensor_rd_data_bits_5_1; // @[Load.scala 97:29:@5751.4]
  assign io_wgt_rd_data_bits_5_2 = tensorLoad_1_io_tensor_rd_data_bits_5_2; // @[Load.scala 97:29:@5752.4]
  assign io_wgt_rd_data_bits_5_3 = tensorLoad_1_io_tensor_rd_data_bits_5_3; // @[Load.scala 97:29:@5753.4]
  assign io_wgt_rd_data_bits_5_4 = tensorLoad_1_io_tensor_rd_data_bits_5_4; // @[Load.scala 97:29:@5754.4]
  assign io_wgt_rd_data_bits_5_5 = tensorLoad_1_io_tensor_rd_data_bits_5_5; // @[Load.scala 97:29:@5755.4]
  assign io_wgt_rd_data_bits_5_6 = tensorLoad_1_io_tensor_rd_data_bits_5_6; // @[Load.scala 97:29:@5756.4]
  assign io_wgt_rd_data_bits_5_7 = tensorLoad_1_io_tensor_rd_data_bits_5_7; // @[Load.scala 97:29:@5757.4]
  assign io_wgt_rd_data_bits_5_8 = tensorLoad_1_io_tensor_rd_data_bits_5_8; // @[Load.scala 97:29:@5758.4]
  assign io_wgt_rd_data_bits_5_9 = tensorLoad_1_io_tensor_rd_data_bits_5_9; // @[Load.scala 97:29:@5759.4]
  assign io_wgt_rd_data_bits_5_10 = tensorLoad_1_io_tensor_rd_data_bits_5_10; // @[Load.scala 97:29:@5760.4]
  assign io_wgt_rd_data_bits_5_11 = tensorLoad_1_io_tensor_rd_data_bits_5_11; // @[Load.scala 97:29:@5761.4]
  assign io_wgt_rd_data_bits_5_12 = tensorLoad_1_io_tensor_rd_data_bits_5_12; // @[Load.scala 97:29:@5762.4]
  assign io_wgt_rd_data_bits_5_13 = tensorLoad_1_io_tensor_rd_data_bits_5_13; // @[Load.scala 97:29:@5763.4]
  assign io_wgt_rd_data_bits_5_14 = tensorLoad_1_io_tensor_rd_data_bits_5_14; // @[Load.scala 97:29:@5764.4]
  assign io_wgt_rd_data_bits_5_15 = tensorLoad_1_io_tensor_rd_data_bits_5_15; // @[Load.scala 97:29:@5765.4]
  assign io_wgt_rd_data_bits_6_0 = tensorLoad_1_io_tensor_rd_data_bits_6_0; // @[Load.scala 97:29:@5766.4]
  assign io_wgt_rd_data_bits_6_1 = tensorLoad_1_io_tensor_rd_data_bits_6_1; // @[Load.scala 97:29:@5767.4]
  assign io_wgt_rd_data_bits_6_2 = tensorLoad_1_io_tensor_rd_data_bits_6_2; // @[Load.scala 97:29:@5768.4]
  assign io_wgt_rd_data_bits_6_3 = tensorLoad_1_io_tensor_rd_data_bits_6_3; // @[Load.scala 97:29:@5769.4]
  assign io_wgt_rd_data_bits_6_4 = tensorLoad_1_io_tensor_rd_data_bits_6_4; // @[Load.scala 97:29:@5770.4]
  assign io_wgt_rd_data_bits_6_5 = tensorLoad_1_io_tensor_rd_data_bits_6_5; // @[Load.scala 97:29:@5771.4]
  assign io_wgt_rd_data_bits_6_6 = tensorLoad_1_io_tensor_rd_data_bits_6_6; // @[Load.scala 97:29:@5772.4]
  assign io_wgt_rd_data_bits_6_7 = tensorLoad_1_io_tensor_rd_data_bits_6_7; // @[Load.scala 97:29:@5773.4]
  assign io_wgt_rd_data_bits_6_8 = tensorLoad_1_io_tensor_rd_data_bits_6_8; // @[Load.scala 97:29:@5774.4]
  assign io_wgt_rd_data_bits_6_9 = tensorLoad_1_io_tensor_rd_data_bits_6_9; // @[Load.scala 97:29:@5775.4]
  assign io_wgt_rd_data_bits_6_10 = tensorLoad_1_io_tensor_rd_data_bits_6_10; // @[Load.scala 97:29:@5776.4]
  assign io_wgt_rd_data_bits_6_11 = tensorLoad_1_io_tensor_rd_data_bits_6_11; // @[Load.scala 97:29:@5777.4]
  assign io_wgt_rd_data_bits_6_12 = tensorLoad_1_io_tensor_rd_data_bits_6_12; // @[Load.scala 97:29:@5778.4]
  assign io_wgt_rd_data_bits_6_13 = tensorLoad_1_io_tensor_rd_data_bits_6_13; // @[Load.scala 97:29:@5779.4]
  assign io_wgt_rd_data_bits_6_14 = tensorLoad_1_io_tensor_rd_data_bits_6_14; // @[Load.scala 97:29:@5780.4]
  assign io_wgt_rd_data_bits_6_15 = tensorLoad_1_io_tensor_rd_data_bits_6_15; // @[Load.scala 97:29:@5781.4]
  assign io_wgt_rd_data_bits_7_0 = tensorLoad_1_io_tensor_rd_data_bits_7_0; // @[Load.scala 97:29:@5782.4]
  assign io_wgt_rd_data_bits_7_1 = tensorLoad_1_io_tensor_rd_data_bits_7_1; // @[Load.scala 97:29:@5783.4]
  assign io_wgt_rd_data_bits_7_2 = tensorLoad_1_io_tensor_rd_data_bits_7_2; // @[Load.scala 97:29:@5784.4]
  assign io_wgt_rd_data_bits_7_3 = tensorLoad_1_io_tensor_rd_data_bits_7_3; // @[Load.scala 97:29:@5785.4]
  assign io_wgt_rd_data_bits_7_4 = tensorLoad_1_io_tensor_rd_data_bits_7_4; // @[Load.scala 97:29:@5786.4]
  assign io_wgt_rd_data_bits_7_5 = tensorLoad_1_io_tensor_rd_data_bits_7_5; // @[Load.scala 97:29:@5787.4]
  assign io_wgt_rd_data_bits_7_6 = tensorLoad_1_io_tensor_rd_data_bits_7_6; // @[Load.scala 97:29:@5788.4]
  assign io_wgt_rd_data_bits_7_7 = tensorLoad_1_io_tensor_rd_data_bits_7_7; // @[Load.scala 97:29:@5789.4]
  assign io_wgt_rd_data_bits_7_8 = tensorLoad_1_io_tensor_rd_data_bits_7_8; // @[Load.scala 97:29:@5790.4]
  assign io_wgt_rd_data_bits_7_9 = tensorLoad_1_io_tensor_rd_data_bits_7_9; // @[Load.scala 97:29:@5791.4]
  assign io_wgt_rd_data_bits_7_10 = tensorLoad_1_io_tensor_rd_data_bits_7_10; // @[Load.scala 97:29:@5792.4]
  assign io_wgt_rd_data_bits_7_11 = tensorLoad_1_io_tensor_rd_data_bits_7_11; // @[Load.scala 97:29:@5793.4]
  assign io_wgt_rd_data_bits_7_12 = tensorLoad_1_io_tensor_rd_data_bits_7_12; // @[Load.scala 97:29:@5794.4]
  assign io_wgt_rd_data_bits_7_13 = tensorLoad_1_io_tensor_rd_data_bits_7_13; // @[Load.scala 97:29:@5795.4]
  assign io_wgt_rd_data_bits_7_14 = tensorLoad_1_io_tensor_rd_data_bits_7_14; // @[Load.scala 97:29:@5796.4]
  assign io_wgt_rd_data_bits_7_15 = tensorLoad_1_io_tensor_rd_data_bits_7_15; // @[Load.scala 97:29:@5797.4]
  assign io_wgt_rd_data_bits_8_0 = tensorLoad_1_io_tensor_rd_data_bits_8_0; // @[Load.scala 97:29:@5798.4]
  assign io_wgt_rd_data_bits_8_1 = tensorLoad_1_io_tensor_rd_data_bits_8_1; // @[Load.scala 97:29:@5799.4]
  assign io_wgt_rd_data_bits_8_2 = tensorLoad_1_io_tensor_rd_data_bits_8_2; // @[Load.scala 97:29:@5800.4]
  assign io_wgt_rd_data_bits_8_3 = tensorLoad_1_io_tensor_rd_data_bits_8_3; // @[Load.scala 97:29:@5801.4]
  assign io_wgt_rd_data_bits_8_4 = tensorLoad_1_io_tensor_rd_data_bits_8_4; // @[Load.scala 97:29:@5802.4]
  assign io_wgt_rd_data_bits_8_5 = tensorLoad_1_io_tensor_rd_data_bits_8_5; // @[Load.scala 97:29:@5803.4]
  assign io_wgt_rd_data_bits_8_6 = tensorLoad_1_io_tensor_rd_data_bits_8_6; // @[Load.scala 97:29:@5804.4]
  assign io_wgt_rd_data_bits_8_7 = tensorLoad_1_io_tensor_rd_data_bits_8_7; // @[Load.scala 97:29:@5805.4]
  assign io_wgt_rd_data_bits_8_8 = tensorLoad_1_io_tensor_rd_data_bits_8_8; // @[Load.scala 97:29:@5806.4]
  assign io_wgt_rd_data_bits_8_9 = tensorLoad_1_io_tensor_rd_data_bits_8_9; // @[Load.scala 97:29:@5807.4]
  assign io_wgt_rd_data_bits_8_10 = tensorLoad_1_io_tensor_rd_data_bits_8_10; // @[Load.scala 97:29:@5808.4]
  assign io_wgt_rd_data_bits_8_11 = tensorLoad_1_io_tensor_rd_data_bits_8_11; // @[Load.scala 97:29:@5809.4]
  assign io_wgt_rd_data_bits_8_12 = tensorLoad_1_io_tensor_rd_data_bits_8_12; // @[Load.scala 97:29:@5810.4]
  assign io_wgt_rd_data_bits_8_13 = tensorLoad_1_io_tensor_rd_data_bits_8_13; // @[Load.scala 97:29:@5811.4]
  assign io_wgt_rd_data_bits_8_14 = tensorLoad_1_io_tensor_rd_data_bits_8_14; // @[Load.scala 97:29:@5812.4]
  assign io_wgt_rd_data_bits_8_15 = tensorLoad_1_io_tensor_rd_data_bits_8_15; // @[Load.scala 97:29:@5813.4]
  assign io_wgt_rd_data_bits_9_0 = tensorLoad_1_io_tensor_rd_data_bits_9_0; // @[Load.scala 97:29:@5814.4]
  assign io_wgt_rd_data_bits_9_1 = tensorLoad_1_io_tensor_rd_data_bits_9_1; // @[Load.scala 97:29:@5815.4]
  assign io_wgt_rd_data_bits_9_2 = tensorLoad_1_io_tensor_rd_data_bits_9_2; // @[Load.scala 97:29:@5816.4]
  assign io_wgt_rd_data_bits_9_3 = tensorLoad_1_io_tensor_rd_data_bits_9_3; // @[Load.scala 97:29:@5817.4]
  assign io_wgt_rd_data_bits_9_4 = tensorLoad_1_io_tensor_rd_data_bits_9_4; // @[Load.scala 97:29:@5818.4]
  assign io_wgt_rd_data_bits_9_5 = tensorLoad_1_io_tensor_rd_data_bits_9_5; // @[Load.scala 97:29:@5819.4]
  assign io_wgt_rd_data_bits_9_6 = tensorLoad_1_io_tensor_rd_data_bits_9_6; // @[Load.scala 97:29:@5820.4]
  assign io_wgt_rd_data_bits_9_7 = tensorLoad_1_io_tensor_rd_data_bits_9_7; // @[Load.scala 97:29:@5821.4]
  assign io_wgt_rd_data_bits_9_8 = tensorLoad_1_io_tensor_rd_data_bits_9_8; // @[Load.scala 97:29:@5822.4]
  assign io_wgt_rd_data_bits_9_9 = tensorLoad_1_io_tensor_rd_data_bits_9_9; // @[Load.scala 97:29:@5823.4]
  assign io_wgt_rd_data_bits_9_10 = tensorLoad_1_io_tensor_rd_data_bits_9_10; // @[Load.scala 97:29:@5824.4]
  assign io_wgt_rd_data_bits_9_11 = tensorLoad_1_io_tensor_rd_data_bits_9_11; // @[Load.scala 97:29:@5825.4]
  assign io_wgt_rd_data_bits_9_12 = tensorLoad_1_io_tensor_rd_data_bits_9_12; // @[Load.scala 97:29:@5826.4]
  assign io_wgt_rd_data_bits_9_13 = tensorLoad_1_io_tensor_rd_data_bits_9_13; // @[Load.scala 97:29:@5827.4]
  assign io_wgt_rd_data_bits_9_14 = tensorLoad_1_io_tensor_rd_data_bits_9_14; // @[Load.scala 97:29:@5828.4]
  assign io_wgt_rd_data_bits_9_15 = tensorLoad_1_io_tensor_rd_data_bits_9_15; // @[Load.scala 97:29:@5829.4]
  assign io_wgt_rd_data_bits_10_0 = tensorLoad_1_io_tensor_rd_data_bits_10_0; // @[Load.scala 97:29:@5830.4]
  assign io_wgt_rd_data_bits_10_1 = tensorLoad_1_io_tensor_rd_data_bits_10_1; // @[Load.scala 97:29:@5831.4]
  assign io_wgt_rd_data_bits_10_2 = tensorLoad_1_io_tensor_rd_data_bits_10_2; // @[Load.scala 97:29:@5832.4]
  assign io_wgt_rd_data_bits_10_3 = tensorLoad_1_io_tensor_rd_data_bits_10_3; // @[Load.scala 97:29:@5833.4]
  assign io_wgt_rd_data_bits_10_4 = tensorLoad_1_io_tensor_rd_data_bits_10_4; // @[Load.scala 97:29:@5834.4]
  assign io_wgt_rd_data_bits_10_5 = tensorLoad_1_io_tensor_rd_data_bits_10_5; // @[Load.scala 97:29:@5835.4]
  assign io_wgt_rd_data_bits_10_6 = tensorLoad_1_io_tensor_rd_data_bits_10_6; // @[Load.scala 97:29:@5836.4]
  assign io_wgt_rd_data_bits_10_7 = tensorLoad_1_io_tensor_rd_data_bits_10_7; // @[Load.scala 97:29:@5837.4]
  assign io_wgt_rd_data_bits_10_8 = tensorLoad_1_io_tensor_rd_data_bits_10_8; // @[Load.scala 97:29:@5838.4]
  assign io_wgt_rd_data_bits_10_9 = tensorLoad_1_io_tensor_rd_data_bits_10_9; // @[Load.scala 97:29:@5839.4]
  assign io_wgt_rd_data_bits_10_10 = tensorLoad_1_io_tensor_rd_data_bits_10_10; // @[Load.scala 97:29:@5840.4]
  assign io_wgt_rd_data_bits_10_11 = tensorLoad_1_io_tensor_rd_data_bits_10_11; // @[Load.scala 97:29:@5841.4]
  assign io_wgt_rd_data_bits_10_12 = tensorLoad_1_io_tensor_rd_data_bits_10_12; // @[Load.scala 97:29:@5842.4]
  assign io_wgt_rd_data_bits_10_13 = tensorLoad_1_io_tensor_rd_data_bits_10_13; // @[Load.scala 97:29:@5843.4]
  assign io_wgt_rd_data_bits_10_14 = tensorLoad_1_io_tensor_rd_data_bits_10_14; // @[Load.scala 97:29:@5844.4]
  assign io_wgt_rd_data_bits_10_15 = tensorLoad_1_io_tensor_rd_data_bits_10_15; // @[Load.scala 97:29:@5845.4]
  assign io_wgt_rd_data_bits_11_0 = tensorLoad_1_io_tensor_rd_data_bits_11_0; // @[Load.scala 97:29:@5846.4]
  assign io_wgt_rd_data_bits_11_1 = tensorLoad_1_io_tensor_rd_data_bits_11_1; // @[Load.scala 97:29:@5847.4]
  assign io_wgt_rd_data_bits_11_2 = tensorLoad_1_io_tensor_rd_data_bits_11_2; // @[Load.scala 97:29:@5848.4]
  assign io_wgt_rd_data_bits_11_3 = tensorLoad_1_io_tensor_rd_data_bits_11_3; // @[Load.scala 97:29:@5849.4]
  assign io_wgt_rd_data_bits_11_4 = tensorLoad_1_io_tensor_rd_data_bits_11_4; // @[Load.scala 97:29:@5850.4]
  assign io_wgt_rd_data_bits_11_5 = tensorLoad_1_io_tensor_rd_data_bits_11_5; // @[Load.scala 97:29:@5851.4]
  assign io_wgt_rd_data_bits_11_6 = tensorLoad_1_io_tensor_rd_data_bits_11_6; // @[Load.scala 97:29:@5852.4]
  assign io_wgt_rd_data_bits_11_7 = tensorLoad_1_io_tensor_rd_data_bits_11_7; // @[Load.scala 97:29:@5853.4]
  assign io_wgt_rd_data_bits_11_8 = tensorLoad_1_io_tensor_rd_data_bits_11_8; // @[Load.scala 97:29:@5854.4]
  assign io_wgt_rd_data_bits_11_9 = tensorLoad_1_io_tensor_rd_data_bits_11_9; // @[Load.scala 97:29:@5855.4]
  assign io_wgt_rd_data_bits_11_10 = tensorLoad_1_io_tensor_rd_data_bits_11_10; // @[Load.scala 97:29:@5856.4]
  assign io_wgt_rd_data_bits_11_11 = tensorLoad_1_io_tensor_rd_data_bits_11_11; // @[Load.scala 97:29:@5857.4]
  assign io_wgt_rd_data_bits_11_12 = tensorLoad_1_io_tensor_rd_data_bits_11_12; // @[Load.scala 97:29:@5858.4]
  assign io_wgt_rd_data_bits_11_13 = tensorLoad_1_io_tensor_rd_data_bits_11_13; // @[Load.scala 97:29:@5859.4]
  assign io_wgt_rd_data_bits_11_14 = tensorLoad_1_io_tensor_rd_data_bits_11_14; // @[Load.scala 97:29:@5860.4]
  assign io_wgt_rd_data_bits_11_15 = tensorLoad_1_io_tensor_rd_data_bits_11_15; // @[Load.scala 97:29:@5861.4]
  assign io_wgt_rd_data_bits_12_0 = tensorLoad_1_io_tensor_rd_data_bits_12_0; // @[Load.scala 97:29:@5862.4]
  assign io_wgt_rd_data_bits_12_1 = tensorLoad_1_io_tensor_rd_data_bits_12_1; // @[Load.scala 97:29:@5863.4]
  assign io_wgt_rd_data_bits_12_2 = tensorLoad_1_io_tensor_rd_data_bits_12_2; // @[Load.scala 97:29:@5864.4]
  assign io_wgt_rd_data_bits_12_3 = tensorLoad_1_io_tensor_rd_data_bits_12_3; // @[Load.scala 97:29:@5865.4]
  assign io_wgt_rd_data_bits_12_4 = tensorLoad_1_io_tensor_rd_data_bits_12_4; // @[Load.scala 97:29:@5866.4]
  assign io_wgt_rd_data_bits_12_5 = tensorLoad_1_io_tensor_rd_data_bits_12_5; // @[Load.scala 97:29:@5867.4]
  assign io_wgt_rd_data_bits_12_6 = tensorLoad_1_io_tensor_rd_data_bits_12_6; // @[Load.scala 97:29:@5868.4]
  assign io_wgt_rd_data_bits_12_7 = tensorLoad_1_io_tensor_rd_data_bits_12_7; // @[Load.scala 97:29:@5869.4]
  assign io_wgt_rd_data_bits_12_8 = tensorLoad_1_io_tensor_rd_data_bits_12_8; // @[Load.scala 97:29:@5870.4]
  assign io_wgt_rd_data_bits_12_9 = tensorLoad_1_io_tensor_rd_data_bits_12_9; // @[Load.scala 97:29:@5871.4]
  assign io_wgt_rd_data_bits_12_10 = tensorLoad_1_io_tensor_rd_data_bits_12_10; // @[Load.scala 97:29:@5872.4]
  assign io_wgt_rd_data_bits_12_11 = tensorLoad_1_io_tensor_rd_data_bits_12_11; // @[Load.scala 97:29:@5873.4]
  assign io_wgt_rd_data_bits_12_12 = tensorLoad_1_io_tensor_rd_data_bits_12_12; // @[Load.scala 97:29:@5874.4]
  assign io_wgt_rd_data_bits_12_13 = tensorLoad_1_io_tensor_rd_data_bits_12_13; // @[Load.scala 97:29:@5875.4]
  assign io_wgt_rd_data_bits_12_14 = tensorLoad_1_io_tensor_rd_data_bits_12_14; // @[Load.scala 97:29:@5876.4]
  assign io_wgt_rd_data_bits_12_15 = tensorLoad_1_io_tensor_rd_data_bits_12_15; // @[Load.scala 97:29:@5877.4]
  assign io_wgt_rd_data_bits_13_0 = tensorLoad_1_io_tensor_rd_data_bits_13_0; // @[Load.scala 97:29:@5878.4]
  assign io_wgt_rd_data_bits_13_1 = tensorLoad_1_io_tensor_rd_data_bits_13_1; // @[Load.scala 97:29:@5879.4]
  assign io_wgt_rd_data_bits_13_2 = tensorLoad_1_io_tensor_rd_data_bits_13_2; // @[Load.scala 97:29:@5880.4]
  assign io_wgt_rd_data_bits_13_3 = tensorLoad_1_io_tensor_rd_data_bits_13_3; // @[Load.scala 97:29:@5881.4]
  assign io_wgt_rd_data_bits_13_4 = tensorLoad_1_io_tensor_rd_data_bits_13_4; // @[Load.scala 97:29:@5882.4]
  assign io_wgt_rd_data_bits_13_5 = tensorLoad_1_io_tensor_rd_data_bits_13_5; // @[Load.scala 97:29:@5883.4]
  assign io_wgt_rd_data_bits_13_6 = tensorLoad_1_io_tensor_rd_data_bits_13_6; // @[Load.scala 97:29:@5884.4]
  assign io_wgt_rd_data_bits_13_7 = tensorLoad_1_io_tensor_rd_data_bits_13_7; // @[Load.scala 97:29:@5885.4]
  assign io_wgt_rd_data_bits_13_8 = tensorLoad_1_io_tensor_rd_data_bits_13_8; // @[Load.scala 97:29:@5886.4]
  assign io_wgt_rd_data_bits_13_9 = tensorLoad_1_io_tensor_rd_data_bits_13_9; // @[Load.scala 97:29:@5887.4]
  assign io_wgt_rd_data_bits_13_10 = tensorLoad_1_io_tensor_rd_data_bits_13_10; // @[Load.scala 97:29:@5888.4]
  assign io_wgt_rd_data_bits_13_11 = tensorLoad_1_io_tensor_rd_data_bits_13_11; // @[Load.scala 97:29:@5889.4]
  assign io_wgt_rd_data_bits_13_12 = tensorLoad_1_io_tensor_rd_data_bits_13_12; // @[Load.scala 97:29:@5890.4]
  assign io_wgt_rd_data_bits_13_13 = tensorLoad_1_io_tensor_rd_data_bits_13_13; // @[Load.scala 97:29:@5891.4]
  assign io_wgt_rd_data_bits_13_14 = tensorLoad_1_io_tensor_rd_data_bits_13_14; // @[Load.scala 97:29:@5892.4]
  assign io_wgt_rd_data_bits_13_15 = tensorLoad_1_io_tensor_rd_data_bits_13_15; // @[Load.scala 97:29:@5893.4]
  assign io_wgt_rd_data_bits_14_0 = tensorLoad_1_io_tensor_rd_data_bits_14_0; // @[Load.scala 97:29:@5894.4]
  assign io_wgt_rd_data_bits_14_1 = tensorLoad_1_io_tensor_rd_data_bits_14_1; // @[Load.scala 97:29:@5895.4]
  assign io_wgt_rd_data_bits_14_2 = tensorLoad_1_io_tensor_rd_data_bits_14_2; // @[Load.scala 97:29:@5896.4]
  assign io_wgt_rd_data_bits_14_3 = tensorLoad_1_io_tensor_rd_data_bits_14_3; // @[Load.scala 97:29:@5897.4]
  assign io_wgt_rd_data_bits_14_4 = tensorLoad_1_io_tensor_rd_data_bits_14_4; // @[Load.scala 97:29:@5898.4]
  assign io_wgt_rd_data_bits_14_5 = tensorLoad_1_io_tensor_rd_data_bits_14_5; // @[Load.scala 97:29:@5899.4]
  assign io_wgt_rd_data_bits_14_6 = tensorLoad_1_io_tensor_rd_data_bits_14_6; // @[Load.scala 97:29:@5900.4]
  assign io_wgt_rd_data_bits_14_7 = tensorLoad_1_io_tensor_rd_data_bits_14_7; // @[Load.scala 97:29:@5901.4]
  assign io_wgt_rd_data_bits_14_8 = tensorLoad_1_io_tensor_rd_data_bits_14_8; // @[Load.scala 97:29:@5902.4]
  assign io_wgt_rd_data_bits_14_9 = tensorLoad_1_io_tensor_rd_data_bits_14_9; // @[Load.scala 97:29:@5903.4]
  assign io_wgt_rd_data_bits_14_10 = tensorLoad_1_io_tensor_rd_data_bits_14_10; // @[Load.scala 97:29:@5904.4]
  assign io_wgt_rd_data_bits_14_11 = tensorLoad_1_io_tensor_rd_data_bits_14_11; // @[Load.scala 97:29:@5905.4]
  assign io_wgt_rd_data_bits_14_12 = tensorLoad_1_io_tensor_rd_data_bits_14_12; // @[Load.scala 97:29:@5906.4]
  assign io_wgt_rd_data_bits_14_13 = tensorLoad_1_io_tensor_rd_data_bits_14_13; // @[Load.scala 97:29:@5907.4]
  assign io_wgt_rd_data_bits_14_14 = tensorLoad_1_io_tensor_rd_data_bits_14_14; // @[Load.scala 97:29:@5908.4]
  assign io_wgt_rd_data_bits_14_15 = tensorLoad_1_io_tensor_rd_data_bits_14_15; // @[Load.scala 97:29:@5909.4]
  assign io_wgt_rd_data_bits_15_0 = tensorLoad_1_io_tensor_rd_data_bits_15_0; // @[Load.scala 97:29:@5910.4]
  assign io_wgt_rd_data_bits_15_1 = tensorLoad_1_io_tensor_rd_data_bits_15_1; // @[Load.scala 97:29:@5911.4]
  assign io_wgt_rd_data_bits_15_2 = tensorLoad_1_io_tensor_rd_data_bits_15_2; // @[Load.scala 97:29:@5912.4]
  assign io_wgt_rd_data_bits_15_3 = tensorLoad_1_io_tensor_rd_data_bits_15_3; // @[Load.scala 97:29:@5913.4]
  assign io_wgt_rd_data_bits_15_4 = tensorLoad_1_io_tensor_rd_data_bits_15_4; // @[Load.scala 97:29:@5914.4]
  assign io_wgt_rd_data_bits_15_5 = tensorLoad_1_io_tensor_rd_data_bits_15_5; // @[Load.scala 97:29:@5915.4]
  assign io_wgt_rd_data_bits_15_6 = tensorLoad_1_io_tensor_rd_data_bits_15_6; // @[Load.scala 97:29:@5916.4]
  assign io_wgt_rd_data_bits_15_7 = tensorLoad_1_io_tensor_rd_data_bits_15_7; // @[Load.scala 97:29:@5917.4]
  assign io_wgt_rd_data_bits_15_8 = tensorLoad_1_io_tensor_rd_data_bits_15_8; // @[Load.scala 97:29:@5918.4]
  assign io_wgt_rd_data_bits_15_9 = tensorLoad_1_io_tensor_rd_data_bits_15_9; // @[Load.scala 97:29:@5919.4]
  assign io_wgt_rd_data_bits_15_10 = tensorLoad_1_io_tensor_rd_data_bits_15_10; // @[Load.scala 97:29:@5920.4]
  assign io_wgt_rd_data_bits_15_11 = tensorLoad_1_io_tensor_rd_data_bits_15_11; // @[Load.scala 97:29:@5921.4]
  assign io_wgt_rd_data_bits_15_12 = tensorLoad_1_io_tensor_rd_data_bits_15_12; // @[Load.scala 97:29:@5922.4]
  assign io_wgt_rd_data_bits_15_13 = tensorLoad_1_io_tensor_rd_data_bits_15_13; // @[Load.scala 97:29:@5923.4]
  assign io_wgt_rd_data_bits_15_14 = tensorLoad_1_io_tensor_rd_data_bits_15_14; // @[Load.scala 97:29:@5924.4]
  assign io_wgt_rd_data_bits_15_15 = tensorLoad_1_io_tensor_rd_data_bits_15_15; // @[Load.scala 97:29:@5925.4]
  assign s_clock = clock; // @[:@5305.4]
  assign s_reset = reset; // @[:@5306.4]
  assign s_io_spost = io_i_post; // @[Load.scala 102:14:@5936.4]
  assign s_io_swait = dec_io_pop_next & _T_5009; // @[Load.scala 103:14:@5940.4]
  assign inst_q_clock = clock; // @[:@5308.4]
  assign inst_q_reset = reset; // @[:@5309.4]
  assign inst_q_io_enq_valid = io_inst_valid; // @[Load.scala 85:17:@5349.4]
  assign inst_q_io_enq_bits = io_inst_bits; // @[Load.scala 85:17:@5348.4]
  assign inst_q_io_deq_ready = _T_5005 | _T_5006; // @[Load.scala 86:23:@5355.4]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Load.scala 53:15:@5313.4]
  assign tensorLoad_0_clock = clock; // @[:@5315.4]
  assign tensorLoad_0_reset = reset; // @[:@5316.4]
  assign tensorLoad_0_io_start = _T_5009 & dec_io_isInput; // @[Load.scala 94:28:@5359.4]
  assign tensorLoad_0_io_inst = inst_q_io_deq_bits; // @[Load.scala 95:27:@5360.4]
  assign tensorLoad_0_io_baddr = io_inp_baddr; // @[Load.scala 96:28:@5361.4]
  assign tensorLoad_0_io_vme_rd_cmd_ready = io_vme_rd_0_cmd_ready; // @[Load.scala 98:18:@5405.4]
  assign tensorLoad_0_io_vme_rd_data_valid = io_vme_rd_0_data_valid; // @[Load.scala 98:18:@5400.4]
  assign tensorLoad_0_io_vme_rd_data_bits = io_vme_rd_0_data_bits; // @[Load.scala 98:18:@5399.4]
  assign tensorLoad_0_io_tensor_rd_idx_valid = io_inp_rd_idx_valid; // @[Load.scala 97:29:@5398.4]
  assign tensorLoad_0_io_tensor_rd_idx_bits = io_inp_rd_idx_bits; // @[Load.scala 97:29:@5397.4]
  assign tensorLoad_1_clock = clock; // @[:@5318.4]
  assign tensorLoad_1_reset = reset; // @[:@5319.4]
  assign tensorLoad_1_io_start = _T_5009 & dec_io_isWeight; // @[Load.scala 94:28:@5409.4]
  assign tensorLoad_1_io_inst = inst_q_io_deq_bits; // @[Load.scala 95:27:@5410.4]
  assign tensorLoad_1_io_baddr = io_wgt_baddr; // @[Load.scala 96:28:@5411.4]
  assign tensorLoad_1_io_vme_rd_cmd_ready = io_vme_rd_1_cmd_ready; // @[Load.scala 98:18:@5935.4]
  assign tensorLoad_1_io_vme_rd_data_valid = io_vme_rd_1_data_valid; // @[Load.scala 98:18:@5930.4]
  assign tensorLoad_1_io_vme_rd_data_bits = io_vme_rd_1_data_bits; // @[Load.scala 98:18:@5929.4]
  assign tensorLoad_1_io_tensor_rd_idx_valid = io_wgt_rd_idx_valid; // @[Load.scala 97:29:@5928.4]
  assign tensorLoad_1_io_tensor_rd_idx_bits = io_wgt_rd_idx_bits; // @[Load.scala 97:29:@5927.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_5000) begin
        if (start) begin
          if (dec_io_isSync) begin
            state <= 2'h1;
          end else begin
            if (_T_5001) begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_5002) begin
          state <= 2'h0;
        end else begin
          if (_T_5003) begin
            if (done) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module LoadUop( // @[:@6004.2]
  input          clock, // @[:@6005.4]
  input          reset, // @[:@6006.4]
  input          io_start, // @[:@6007.4]
  output         io_done, // @[:@6007.4]
  input  [127:0] io_inst, // @[:@6007.4]
  input  [31:0]  io_baddr, // @[:@6007.4]
  input          io_vme_rd_cmd_ready, // @[:@6007.4]
  output         io_vme_rd_cmd_valid, // @[:@6007.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@6007.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@6007.4]
  output         io_vme_rd_data_ready, // @[:@6007.4]
  input          io_vme_rd_data_valid, // @[:@6007.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@6007.4]
  input          io_uop_idx_valid, // @[:@6007.4]
  input  [10:0]  io_uop_idx_bits, // @[:@6007.4]
  output         io_uop_data_valid, // @[:@6007.4]
  output [9:0]   io_uop_data_bits_u2, // @[:@6007.4]
  output [10:0]  io_uop_data_bits_u1, // @[:@6007.4]
  output [10:0]  io_uop_data_bits_u0 // @[:@6007.4]
);
  reg [31:0] mem_0 [0:1023]; // @[LoadUop.scala 163:24:@6241.4]
  reg [31:0] _RAND_0;
  wire [31:0] mem_0_memRead_data; // @[LoadUop.scala 163:24:@6241.4]
  wire [9:0] mem_0_memRead_addr; // @[LoadUop.scala 163:24:@6241.4]
  wire [31:0] mem_0__T_564_data; // @[LoadUop.scala 163:24:@6241.4]
  wire [9:0] mem_0__T_564_addr; // @[LoadUop.scala 163:24:@6241.4]
  wire  mem_0__T_564_mask; // @[LoadUop.scala 163:24:@6241.4]
  wire  mem_0__T_564_en; // @[LoadUop.scala 163:24:@6241.4]
  reg [31:0] mem_1 [0:1023]; // @[LoadUop.scala 163:24:@6241.4]
  reg [31:0] _RAND_1;
  wire [31:0] mem_1_memRead_data; // @[LoadUop.scala 163:24:@6241.4]
  wire [9:0] mem_1_memRead_addr; // @[LoadUop.scala 163:24:@6241.4]
  wire [31:0] mem_1__T_564_data; // @[LoadUop.scala 163:24:@6241.4]
  wire [9:0] mem_1__T_564_addr; // @[LoadUop.scala 163:24:@6241.4]
  wire  mem_1__T_564_mask; // @[LoadUop.scala 163:24:@6241.4]
  wire  mem_1__T_564_en; // @[LoadUop.scala 163:24:@6241.4]
  wire [15:0] dec_sram_offset; // @[LoadUop.scala 75:29:@6024.4]
  wire [31:0] dec_dram_offset; // @[LoadUop.scala 75:29:@6026.4]
  wire [15:0] dec_xsize; // @[LoadUop.scala 75:29:@6032.4]
  reg [31:0] raddr; // @[LoadUop.scala 76:18:@6044.4]
  reg [31:0] _RAND_2;
  reg [7:0] xcnt; // @[LoadUop.scala 77:17:@6045.4]
  reg [31:0] _RAND_3;
  reg [7:0] xlen; // @[LoadUop.scala 78:17:@6046.4]
  reg [31:0] _RAND_4;
  reg [15:0] xrem; // @[LoadUop.scala 79:17:@6047.4]
  reg [31:0] _RAND_5;
  wire [14:0] _T_67; // @[LoadUop.scala 80:26:@6048.4]
  wire  _T_68; // @[LoadUop.scala 80:58:@6049.4]
  wire [14:0] _GEN_89; // @[LoadUop.scala 80:47:@6050.4]
  wire [15:0] _T_69; // @[LoadUop.scala 80:47:@6050.4]
  wire [14:0] _T_70; // @[LoadUop.scala 80:47:@6051.4]
  wire [15:0] _GEN_6; // @[LoadUop.scala 80:81:@6052.4]
  wire [1:0] _T_72; // @[LoadUop.scala 80:81:@6052.4]
  wire [14:0] _GEN_90; // @[LoadUop.scala 80:62:@6053.4]
  wire [15:0] _T_73; // @[LoadUop.scala 80:62:@6053.4]
  wire [14:0] _T_74; // @[LoadUop.scala 80:62:@6054.4]
  wire [15:0] _T_76; // @[LoadUop.scala 80:88:@6055.4]
  wire [15:0] _T_77; // @[LoadUop.scala 80:88:@6056.4]
  wire [14:0] xsize; // @[LoadUop.scala 80:88:@6057.4]
  wire [31:0] _GEN_31; // @[LoadUop.scala 84:36:@6058.4]
  wire [1:0] _T_79; // @[LoadUop.scala 84:36:@6058.4]
  wire  dram_even; // @[LoadUop.scala 84:43:@6059.4]
  wire  sram_even; // @[LoadUop.scala 85:43:@6061.4]
  wire [15:0] _GEN_36; // @[LoadUop.scala 86:31:@6062.4]
  wire [1:0] _T_85; // @[LoadUop.scala 86:31:@6062.4]
  wire  sizeIsEven; // @[LoadUop.scala 86:38:@6063.4]
  reg [1:0] state; // @[LoadUop.scala 89:22:@6064.4]
  reg [31:0] _RAND_6;
  wire  _T_88; // @[Conditional.scala 37:30:@6065.4]
  wire  _T_89; // @[LoadUop.scala 96:20:@6069.8]
  wire [9:0] _T_92; // @[LoadUop.scala 100:24:@6075.10]
  wire [9:0] _T_93; // @[LoadUop.scala 100:24:@6076.10]
  wire [8:0] _T_94; // @[LoadUop.scala 100:24:@6077.10]
  wire [15:0] _T_95; // @[LoadUop.scala 101:25:@6079.10]
  wire [15:0] _T_96; // @[LoadUop.scala 101:25:@6080.10]
  wire [14:0] _T_97; // @[LoadUop.scala 101:25:@6081.10]
  wire [14:0] _GEN_0; // @[LoadUop.scala 96:28:@6070.8]
  wire [14:0] _GEN_1; // @[LoadUop.scala 96:28:@6070.8]
  wire [1:0] _GEN_2; // @[LoadUop.scala 94:22:@6067.6]
  wire [14:0] _GEN_3; // @[LoadUop.scala 94:22:@6067.6]
  wire [15:0] _GEN_4; // @[LoadUop.scala 94:22:@6067.6]
  wire  _T_98; // @[Conditional.scala 37:30:@6087.6]
  wire [1:0] _GEN_5; // @[LoadUop.scala 106:33:@6089.8]
  wire  _T_99; // @[Conditional.scala 37:30:@6094.8]
  wire  _T_100; // @[LoadUop.scala 112:19:@6097.12]
  wire  _T_102; // @[LoadUop.scala 113:21:@6099.14]
  wire [32:0] _T_103; // @[LoadUop.scala 116:28:@6104.16]
  wire [31:0] _T_104; // @[LoadUop.scala 116:28:@6105.16]
  wire  _T_105; // @[LoadUop.scala 117:23:@6107.16]
  wire [16:0] _T_111; // @[LoadUop.scala 125:28:@6119.18]
  wire [16:0] _T_112; // @[LoadUop.scala 125:28:@6120.18]
  wire [15:0] _T_113; // @[LoadUop.scala 125:28:@6121.18]
  wire [15:0] _GEN_7; // @[LoadUop.scala 117:31:@6108.16]
  wire [15:0] _GEN_8; // @[LoadUop.scala 117:31:@6108.16]
  wire [1:0] _GEN_9; // @[LoadUop.scala 113:30:@6100.14]
  wire [31:0] _GEN_10; // @[LoadUop.scala 113:30:@6100.14]
  wire [15:0] _GEN_11; // @[LoadUop.scala 113:30:@6100.14]
  wire [15:0] _GEN_12; // @[LoadUop.scala 113:30:@6100.14]
  wire [1:0] _GEN_13; // @[LoadUop.scala 112:29:@6098.12]
  wire [31:0] _GEN_14; // @[LoadUop.scala 112:29:@6098.12]
  wire [15:0] _GEN_15; // @[LoadUop.scala 112:29:@6098.12]
  wire [15:0] _GEN_16; // @[LoadUop.scala 112:29:@6098.12]
  wire [1:0] _GEN_17; // @[LoadUop.scala 111:34:@6096.10]
  wire [31:0] _GEN_18; // @[LoadUop.scala 111:34:@6096.10]
  wire [15:0] _GEN_19; // @[LoadUop.scala 111:34:@6096.10]
  wire [15:0] _GEN_20; // @[LoadUop.scala 111:34:@6096.10]
  wire [1:0] _GEN_21; // @[Conditional.scala 39:67:@6095.8]
  wire [31:0] _GEN_22; // @[Conditional.scala 39:67:@6095.8]
  wire [15:0] _GEN_23; // @[Conditional.scala 39:67:@6095.8]
  wire [15:0] _GEN_24; // @[Conditional.scala 39:67:@6095.8]
  wire [1:0] _GEN_25; // @[Conditional.scala 39:67:@6088.6]
  wire [31:0] _GEN_26; // @[Conditional.scala 39:67:@6088.6]
  wire [15:0] _GEN_27; // @[Conditional.scala 39:67:@6088.6]
  wire [15:0] _GEN_28; // @[Conditional.scala 39:67:@6088.6]
  wire [1:0] _GEN_29; // @[Conditional.scala 40:58:@6066.4]
  wire [15:0] _GEN_30; // @[Conditional.scala 40:58:@6066.4]
  wire [31:0] _GEN_32; // @[Conditional.scala 40:58:@6066.4]
  wire  _T_214; // @[LoadUop.scala 135:14:@6192.4]
  wire [33:0] _GEN_91; // @[LoadUop.scala 137:58:@6195.8]
  wire [33:0] _T_215; // @[LoadUop.scala 137:58:@6195.8]
  wire [33:0] _T_216; // @[LoadUop.scala 137:39:@6196.8]
  wire [33:0] _GEN_92; // @[LoadUop.scala 137:25:@6197.8]
  wire [33:0] _T_217; // @[LoadUop.scala 137:25:@6197.8]
  wire [34:0] _T_222; // @[LoadUop.scala 139:84:@6204.8]
  wire [34:0] _T_223; // @[LoadUop.scala 139:84:@6205.8]
  wire [33:0] _T_224; // @[LoadUop.scala 139:84:@6206.8]
  wire [33:0] _GEN_33; // @[LoadUop.scala 136:21:@6194.6]
  wire [33:0] _GEN_34; // @[LoadUop.scala 135:25:@6193.4]
  wire  _T_226; // @[LoadUop.scala 147:33:@6214.4]
  wire  _T_227; // @[LoadUop.scala 149:14:@6216.4]
  wire  _T_229; // @[Decoupled.scala 37:37:@6221.6]
  wire [8:0] _T_231; // @[LoadUop.scala 152:18:@6223.8]
  wire [7:0] _T_232; // @[LoadUop.scala 152:18:@6224.8]
  wire [7:0] _GEN_35; // @[LoadUop.scala 151:37:@6222.6]
  reg [9:0] waddr; // @[LoadUop.scala 155:18:@6227.4]
  reg [31:0] _RAND_7;
  wire [14:0] _T_235; // @[LoadUop.scala 157:30:@6230.6]
  wire [10:0] _T_238; // @[LoadUop.scala 159:20:@6236.8]
  wire [9:0] _T_239; // @[LoadUop.scala 159:20:@6237.8]
  wire [9:0] _GEN_37; // @[LoadUop.scala 158:37:@6235.6]
  wire [14:0] _GEN_38; // @[LoadUop.scala 156:25:@6229.4]
  reg  wmask_0; // @[LoadUop.scala 164:18:@6242.4]
  reg [31:0] _RAND_8;
  reg  wmask_1; // @[LoadUop.scala 164:18:@6242.4]
  reg [31:0] _RAND_9;
  wire  _T_297; // @[Decoupled.scala 37:37:@6256.8]
  wire  _T_299; // @[LoadUop.scala 170:22:@6258.10]
  wire  _GEN_40; // @[LoadUop.scala 170:31:@6259.10]
  wire [8:0] _T_350; // @[LoadUop.scala 176:27:@6285.12]
  wire [8:0] _T_351; // @[LoadUop.scala 176:27:@6286.12]
  wire [7:0] _T_352; // @[LoadUop.scala 176:27:@6287.12]
  wire  _T_353; // @[LoadUop.scala 176:18:@6288.12]
  wire  _T_356; // @[LoadUop.scala 176:34:@6290.12]
  wire  _GEN_42; // @[LoadUop.scala 176:53:@6291.12]
  wire  _GEN_43; // @[LoadUop.scala 175:39:@6284.10]
  wire  _GEN_44; // @[LoadUop.scala 175:39:@6284.10]
  wire  _GEN_45; // @[LoadUop.scala 169:38:@6257.8]
  wire  _GEN_46; // @[LoadUop.scala 169:38:@6257.8]
  wire  _GEN_47; // @[LoadUop.scala 167:22:@6244.6]
  wire  _GEN_48; // @[LoadUop.scala 167:22:@6244.6]
  wire  _T_436; // @[LoadUop.scala 186:23:@6335.10]
  wire  _T_439; // @[LoadUop.scala 186:48:@6337.10]
  wire  _GEN_50; // @[LoadUop.scala 186:67:@6338.10]
  wire  _GEN_52; // @[LoadUop.scala 185:39:@6330.8]
  wire  _GEN_53; // @[LoadUop.scala 183:32:@6317.6]
  wire  _GEN_54; // @[LoadUop.scala 183:32:@6317.6]
  wire [31:0] _T_509; // @[LoadUop.scala 194:40:@6365.4]
  wire [31:0] _T_510; // @[LoadUop.scala 194:40:@6367.4]
  wire  _T_512; // @[LoadUop.scala 195:18:@6371.4]
  wire  _T_513; // @[LoadUop.scala 195:30:@6372.4]
  wire  _T_538; // @[LoadUop.scala 197:24:@6384.6]
  wire  _T_539; // @[LoadUop.scala 197:36:@6385.6]
  wire [31:0] _GEN_57; // @[LoadUop.scala 197:50:@6386.6]
  reg  _T_579; // @[LoadUop.scala 206:31:@6406.4]
  reg [31:0] _RAND_10;
  wire [10:0] _GEN_39; // @[LoadUop.scala 208:30:@6409.4]
  wire [1:0] sIdx; // @[LoadUop.scala 208:30:@6409.4]
  wire [9:0] rIdx; // @[LoadUop.scala 209:30:@6410.4]
  wire  _GEN_72; // @[LoadUop.scala 210:25:@6413.4]
  wire [63:0] _T_599; // @[LoadUop.scala 211:23:@6419.4]
  wire [31:0] sWord_0; // @[LoadUop.scala 211:38:@6423.4]
  wire [31:0] sWord_1; // @[LoadUop.scala 211:38:@6425.4]
  wire  _T_625; // @[:@6427.4]
  wire [31:0] _GEN_76; // @[:@6430.4]
  wire  _T_633; // @[LoadUop.scala 217:34:@6441.4]
  wire  _T_635; // @[LoadUop.scala 217:57:@6443.4]
  reg [9:0] mem_0_memRead_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [9:0] mem_1_memRead_addr_pipe_0;
  reg [31:0] _RAND_12;
  assign mem_0_memRead_addr = mem_0_memRead_addr_pipe_0;
  assign mem_0_memRead_data = mem_0[mem_0_memRead_addr]; // @[LoadUop.scala 163:24:@6241.4]
  assign mem_0__T_564_data = _T_513 ? _T_510 : _T_509;
  assign mem_0__T_564_addr = waddr;
  assign mem_0__T_564_mask = wmask_0;
  assign mem_0__T_564_en = io_vme_rd_data_ready & io_vme_rd_data_valid;
  assign mem_1_memRead_addr = mem_1_memRead_addr_pipe_0;
  assign mem_1_memRead_data = mem_1[mem_1_memRead_addr]; // @[LoadUop.scala 163:24:@6241.4]
  assign mem_1__T_564_data = _T_513 ? _T_510 : _GEN_57;
  assign mem_1__T_564_addr = waddr;
  assign mem_1__T_564_mask = wmask_1;
  assign mem_1__T_564_en = io_vme_rd_data_ready & io_vme_rd_data_valid;
  assign dec_sram_offset = io_inst[24:9]; // @[LoadUop.scala 75:29:@6024.4]
  assign dec_dram_offset = io_inst[56:25]; // @[LoadUop.scala 75:29:@6026.4]
  assign dec_xsize = io_inst[95:80]; // @[LoadUop.scala 75:29:@6032.4]
  assign _T_67 = dec_xsize[15:1]; // @[LoadUop.scala 80:26:@6048.4]
  assign _T_68 = dec_xsize[0]; // @[LoadUop.scala 80:58:@6049.4]
  assign _GEN_89 = {{14'd0}, _T_68}; // @[LoadUop.scala 80:47:@6050.4]
  assign _T_69 = _T_67 + _GEN_89; // @[LoadUop.scala 80:47:@6050.4]
  assign _T_70 = _T_67 + _GEN_89; // @[LoadUop.scala 80:47:@6051.4]
  assign _GEN_6 = dec_sram_offset % 16'h2; // @[LoadUop.scala 80:81:@6052.4]
  assign _T_72 = _GEN_6[1:0]; // @[LoadUop.scala 80:81:@6052.4]
  assign _GEN_90 = {{13'd0}, _T_72}; // @[LoadUop.scala 80:62:@6053.4]
  assign _T_73 = _T_70 + _GEN_90; // @[LoadUop.scala 80:62:@6053.4]
  assign _T_74 = _T_70 + _GEN_90; // @[LoadUop.scala 80:62:@6054.4]
  assign _T_76 = _T_74 - 15'h1; // @[LoadUop.scala 80:88:@6055.4]
  assign _T_77 = $unsigned(_T_76); // @[LoadUop.scala 80:88:@6056.4]
  assign xsize = _T_77[14:0]; // @[LoadUop.scala 80:88:@6057.4]
  assign _GEN_31 = dec_dram_offset % 32'h2; // @[LoadUop.scala 84:36:@6058.4]
  assign _T_79 = _GEN_31[1:0]; // @[LoadUop.scala 84:36:@6058.4]
  assign dram_even = _T_79 == 2'h0; // @[LoadUop.scala 84:43:@6059.4]
  assign sram_even = _T_72 == 2'h0; // @[LoadUop.scala 85:43:@6061.4]
  assign _GEN_36 = dec_xsize % 16'h2; // @[LoadUop.scala 86:31:@6062.4]
  assign _T_85 = _GEN_36[1:0]; // @[LoadUop.scala 86:31:@6062.4]
  assign sizeIsEven = _T_85 == 2'h0; // @[LoadUop.scala 86:38:@6063.4]
  assign _T_88 = 2'h0 == state; // @[Conditional.scala 37:30:@6065.4]
  assign _T_89 = xsize < 15'h100; // @[LoadUop.scala 96:20:@6069.8]
  assign _T_92 = 9'h100 - 9'h1; // @[LoadUop.scala 100:24:@6075.10]
  assign _T_93 = $unsigned(_T_92); // @[LoadUop.scala 100:24:@6076.10]
  assign _T_94 = _T_93[8:0]; // @[LoadUop.scala 100:24:@6077.10]
  assign _T_95 = xsize - 15'h100; // @[LoadUop.scala 101:25:@6079.10]
  assign _T_96 = $unsigned(_T_95); // @[LoadUop.scala 101:25:@6080.10]
  assign _T_97 = _T_96[14:0]; // @[LoadUop.scala 101:25:@6081.10]
  assign _GEN_0 = _T_89 ? xsize : {{6'd0}, _T_94}; // @[LoadUop.scala 96:28:@6070.8]
  assign _GEN_1 = _T_89 ? 15'h0 : _T_97; // @[LoadUop.scala 96:28:@6070.8]
  assign _GEN_2 = io_start ? 2'h1 : state; // @[LoadUop.scala 94:22:@6067.6]
  assign _GEN_3 = io_start ? _GEN_0 : {{7'd0}, xlen}; // @[LoadUop.scala 94:22:@6067.6]
  assign _GEN_4 = io_start ? {{1'd0}, _GEN_1} : xrem; // @[LoadUop.scala 94:22:@6067.6]
  assign _T_98 = 2'h1 == state; // @[Conditional.scala 37:30:@6087.6]
  assign _GEN_5 = io_vme_rd_cmd_ready ? 2'h2 : state; // @[LoadUop.scala 106:33:@6089.8]
  assign _T_99 = 2'h2 == state; // @[Conditional.scala 37:30:@6094.8]
  assign _T_100 = xcnt == xlen; // @[LoadUop.scala 112:19:@6097.12]
  assign _T_102 = xrem == 16'h0; // @[LoadUop.scala 113:21:@6099.14]
  assign _T_103 = raddr + 32'h800; // @[LoadUop.scala 116:28:@6104.16]
  assign _T_104 = raddr + 32'h800; // @[LoadUop.scala 116:28:@6105.16]
  assign _T_105 = xrem < 16'h100; // @[LoadUop.scala 117:23:@6107.16]
  assign _T_111 = xrem - 16'h100; // @[LoadUop.scala 125:28:@6119.18]
  assign _T_112 = $unsigned(_T_111); // @[LoadUop.scala 125:28:@6120.18]
  assign _T_113 = _T_112[15:0]; // @[LoadUop.scala 125:28:@6121.18]
  assign _GEN_7 = _T_105 ? xrem : {{7'd0}, _T_94}; // @[LoadUop.scala 117:31:@6108.16]
  assign _GEN_8 = _T_105 ? 16'h0 : _T_113; // @[LoadUop.scala 117:31:@6108.16]
  assign _GEN_9 = _T_102 ? 2'h0 : 2'h1; // @[LoadUop.scala 113:30:@6100.14]
  assign _GEN_10 = _T_102 ? raddr : _T_104; // @[LoadUop.scala 113:30:@6100.14]
  assign _GEN_11 = _T_102 ? {{8'd0}, xlen} : _GEN_7; // @[LoadUop.scala 113:30:@6100.14]
  assign _GEN_12 = _T_102 ? xrem : _GEN_8; // @[LoadUop.scala 113:30:@6100.14]
  assign _GEN_13 = _T_100 ? _GEN_9 : state; // @[LoadUop.scala 112:29:@6098.12]
  assign _GEN_14 = _T_100 ? _GEN_10 : raddr; // @[LoadUop.scala 112:29:@6098.12]
  assign _GEN_15 = _T_100 ? _GEN_11 : {{8'd0}, xlen}; // @[LoadUop.scala 112:29:@6098.12]
  assign _GEN_16 = _T_100 ? _GEN_12 : xrem; // @[LoadUop.scala 112:29:@6098.12]
  assign _GEN_17 = io_vme_rd_data_valid ? _GEN_13 : state; // @[LoadUop.scala 111:34:@6096.10]
  assign _GEN_18 = io_vme_rd_data_valid ? _GEN_14 : raddr; // @[LoadUop.scala 111:34:@6096.10]
  assign _GEN_19 = io_vme_rd_data_valid ? _GEN_15 : {{8'd0}, xlen}; // @[LoadUop.scala 111:34:@6096.10]
  assign _GEN_20 = io_vme_rd_data_valid ? _GEN_16 : xrem; // @[LoadUop.scala 111:34:@6096.10]
  assign _GEN_21 = _T_99 ? _GEN_17 : state; // @[Conditional.scala 39:67:@6095.8]
  assign _GEN_22 = _T_99 ? _GEN_18 : raddr; // @[Conditional.scala 39:67:@6095.8]
  assign _GEN_23 = _T_99 ? _GEN_19 : {{8'd0}, xlen}; // @[Conditional.scala 39:67:@6095.8]
  assign _GEN_24 = _T_99 ? _GEN_20 : xrem; // @[Conditional.scala 39:67:@6095.8]
  assign _GEN_25 = _T_98 ? _GEN_5 : _GEN_21; // @[Conditional.scala 39:67:@6088.6]
  assign _GEN_26 = _T_98 ? raddr : _GEN_22; // @[Conditional.scala 39:67:@6088.6]
  assign _GEN_27 = _T_98 ? {{8'd0}, xlen} : _GEN_23; // @[Conditional.scala 39:67:@6088.6]
  assign _GEN_28 = _T_98 ? xrem : _GEN_24; // @[Conditional.scala 39:67:@6088.6]
  assign _GEN_29 = _T_88 ? _GEN_2 : _GEN_25; // @[Conditional.scala 40:58:@6066.4]
  assign _GEN_30 = _T_88 ? {{1'd0}, _GEN_3} : _GEN_27; // @[Conditional.scala 40:58:@6066.4]
  assign _GEN_32 = _T_88 ? raddr : _GEN_26; // @[Conditional.scala 40:58:@6066.4]
  assign _T_214 = state == 2'h0; // @[LoadUop.scala 135:14:@6192.4]
  assign _GEN_91 = {{2'd0}, dec_dram_offset}; // @[LoadUop.scala 137:58:@6195.8]
  assign _T_215 = _GEN_91 << 2; // @[LoadUop.scala 137:58:@6195.8]
  assign _T_216 = 34'hffffffff & _T_215; // @[LoadUop.scala 137:39:@6196.8]
  assign _GEN_92 = {{2'd0}, io_baddr}; // @[LoadUop.scala 137:25:@6197.8]
  assign _T_217 = _GEN_92 | _T_216; // @[LoadUop.scala 137:25:@6197.8]
  assign _T_222 = _T_217 - 34'h4; // @[LoadUop.scala 139:84:@6204.8]
  assign _T_223 = $unsigned(_T_222); // @[LoadUop.scala 139:84:@6205.8]
  assign _T_224 = _T_223[33:0]; // @[LoadUop.scala 139:84:@6206.8]
  assign _GEN_33 = dram_even ? _T_217 : _T_224; // @[LoadUop.scala 136:21:@6194.6]
  assign _GEN_34 = _T_214 ? _GEN_33 : {{2'd0}, _GEN_32}; // @[LoadUop.scala 135:25:@6193.4]
  assign _T_226 = state == 2'h2; // @[LoadUop.scala 147:33:@6214.4]
  assign _T_227 = state != 2'h2; // @[LoadUop.scala 149:14:@6216.4]
  assign _T_229 = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[Decoupled.scala 37:37:@6221.6]
  assign _T_231 = xcnt + 8'h1; // @[LoadUop.scala 152:18:@6223.8]
  assign _T_232 = xcnt + 8'h1; // @[LoadUop.scala 152:18:@6224.8]
  assign _GEN_35 = _T_229 ? _T_232 : xcnt; // @[LoadUop.scala 151:37:@6222.6]
  assign _T_235 = dec_sram_offset[15:1]; // @[LoadUop.scala 157:30:@6230.6]
  assign _T_238 = waddr + 10'h1; // @[LoadUop.scala 159:20:@6236.8]
  assign _T_239 = waddr + 10'h1; // @[LoadUop.scala 159:20:@6237.8]
  assign _GEN_37 = _T_229 ? _T_239 : waddr; // @[LoadUop.scala 158:37:@6235.6]
  assign _GEN_38 = _T_214 ? _T_235 : {{5'd0}, _GEN_37}; // @[LoadUop.scala 156:25:@6229.4]
  assign _T_297 = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[Decoupled.scala 37:37:@6256.8]
  assign _T_299 = dec_xsize == 16'h1; // @[LoadUop.scala 170:22:@6258.10]
  assign _GEN_40 = _T_299 ? 1'h0 : 1'h1; // @[LoadUop.scala 170:31:@6259.10]
  assign _T_350 = xlen - 8'h1; // @[LoadUop.scala 176:27:@6285.12]
  assign _T_351 = $unsigned(_T_350); // @[LoadUop.scala 176:27:@6286.12]
  assign _T_352 = _T_351[7:0]; // @[LoadUop.scala 176:27:@6287.12]
  assign _T_353 = xcnt == _T_352; // @[LoadUop.scala 176:18:@6288.12]
  assign _T_356 = _T_353 & _T_102; // @[LoadUop.scala 176:34:@6290.12]
  assign _GEN_42 = _T_356 ? 1'h0 : 1'h1; // @[LoadUop.scala 176:53:@6291.12]
  assign _GEN_43 = _T_229 ? 1'h1 : wmask_0; // @[LoadUop.scala 175:39:@6284.10]
  assign _GEN_44 = _T_229 ? _GEN_42 : wmask_1; // @[LoadUop.scala 175:39:@6284.10]
  assign _GEN_45 = _T_297 ? 1'h1 : _GEN_43; // @[LoadUop.scala 169:38:@6257.8]
  assign _GEN_46 = _T_297 ? _GEN_40 : _GEN_44; // @[LoadUop.scala 169:38:@6257.8]
  assign _GEN_47 = sizeIsEven ? 1'h1 : _GEN_45; // @[LoadUop.scala 167:22:@6244.6]
  assign _GEN_48 = sizeIsEven ? 1'h1 : _GEN_46; // @[LoadUop.scala 167:22:@6244.6]
  assign _T_436 = sizeIsEven & _T_353; // @[LoadUop.scala 186:23:@6335.10]
  assign _T_439 = _T_436 & _T_102; // @[LoadUop.scala 186:48:@6337.10]
  assign _GEN_50 = _T_439 ? 1'h0 : 1'h1; // @[LoadUop.scala 186:67:@6338.10]
  assign _GEN_52 = _T_229 ? _GEN_50 : wmask_1; // @[LoadUop.scala 185:39:@6330.8]
  assign _GEN_53 = _T_297 ? 1'h0 : _GEN_43; // @[LoadUop.scala 183:32:@6317.6]
  assign _GEN_54 = _T_297 ? 1'h1 : _GEN_52; // @[LoadUop.scala 183:32:@6317.6]
  assign _T_509 = io_vme_rd_data_bits[31:0]; // @[LoadUop.scala 194:40:@6365.4]
  assign _T_510 = io_vme_rd_data_bits[63:32]; // @[LoadUop.scala 194:40:@6367.4]
  assign _T_512 = dram_even == 1'h0; // @[LoadUop.scala 195:18:@6371.4]
  assign _T_513 = _T_512 & sram_even; // @[LoadUop.scala 195:30:@6372.4]
  assign _T_538 = sram_even == 1'h0; // @[LoadUop.scala 197:24:@6384.6]
  assign _T_539 = _T_538 & dram_even; // @[LoadUop.scala 197:36:@6385.6]
  assign _GEN_57 = _T_539 ? _T_509 : _T_510; // @[LoadUop.scala 197:50:@6386.6]
  assign _GEN_39 = io_uop_idx_bits % 11'h2; // @[LoadUop.scala 208:30:@6409.4]
  assign sIdx = _GEN_39[1:0]; // @[LoadUop.scala 208:30:@6409.4]
  assign rIdx = io_uop_idx_bits[10:1]; // @[LoadUop.scala 209:30:@6410.4]
  assign _GEN_72 = io_uop_idx_valid; // @[LoadUop.scala 210:25:@6413.4]
  assign _T_599 = {mem_1_memRead_data,mem_0_memRead_data}; // @[LoadUop.scala 211:23:@6419.4]
  assign sWord_0 = _T_599[31:0]; // @[LoadUop.scala 211:38:@6423.4]
  assign sWord_1 = _T_599[63:32]; // @[LoadUop.scala 211:38:@6425.4]
  assign _T_625 = sIdx[0]; // @[:@6427.4]
  assign _GEN_76 = _T_625 ? sWord_1 : sWord_0; // @[:@6430.4]
  assign _T_633 = _T_226 & io_vme_rd_data_valid; // @[LoadUop.scala 217:34:@6441.4]
  assign _T_635 = _T_633 & _T_100; // @[LoadUop.scala 217:57:@6443.4]
  assign io_done = _T_635 & _T_102; // @[LoadUop.scala 217:11:@6446.4]
  assign io_vme_rd_cmd_valid = state == 2'h1; // @[LoadUop.scala 143:23:@6211.4]
  assign io_vme_rd_cmd_bits_addr = raddr; // @[LoadUop.scala 144:27:@6212.4]
  assign io_vme_rd_cmd_bits_len = xlen; // @[LoadUop.scala 145:26:@6213.4]
  assign io_vme_rd_data_ready = state == 2'h2; // @[LoadUop.scala 147:24:@6215.4]
  assign io_uop_data_valid = _T_579; // @[LoadUop.scala 206:21:@6408.4]
  assign io_uop_data_bits_u2 = _GEN_76[31:22]; // @[LoadUop.scala 214:20:@6439.4]
  assign io_uop_data_bits_u1 = _GEN_76[21:11]; // @[LoadUop.scala 214:20:@6438.4]
  assign io_uop_data_bits_u0 = _GEN_76[10:0]; // @[LoadUop.scala 214:20:@6437.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem_0[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem_1[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  raddr = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  xcnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xlen = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  xrem = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  waddr = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wmask_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wmask_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_579 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_0_memRead_addr_pipe_0 = _RAND_11[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mem_1_memRead_addr_pipe_0 = _RAND_12[9:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem_0__T_564_en & mem_0__T_564_mask) begin
      mem_0[mem_0__T_564_addr] <= mem_0__T_564_data; // @[LoadUop.scala 163:24:@6241.4]
    end
    if(mem_1__T_564_en & mem_1__T_564_mask) begin
      mem_1[mem_1__T_564_addr] <= mem_1__T_564_data; // @[LoadUop.scala 163:24:@6241.4]
    end
    raddr <= _GEN_34[31:0];
    if (_T_227) begin
      xcnt <= 8'h0;
    end else begin
      if (_T_229) begin
        xcnt <= _T_232;
      end
    end
    xlen <= _GEN_30[7:0];
    if (_T_88) begin
      if (io_start) begin
        xrem <= {{1'd0}, _GEN_1};
      end
    end else begin
      if (!(_T_98)) begin
        if (_T_99) begin
          if (io_vme_rd_data_valid) begin
            if (_T_100) begin
              if (!(_T_102)) begin
                if (_T_105) begin
                  xrem <= 16'h0;
                end else begin
                  xrem <= _T_113;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_88) begin
        if (io_start) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_98) begin
          if (io_vme_rd_cmd_ready) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_99) begin
            if (io_vme_rd_data_valid) begin
              if (_T_100) begin
                if (_T_102) begin
                  state <= 2'h0;
                end else begin
                  state <= 2'h1;
                end
              end
            end
          end
        end
      end
    end
    waddr <= _GEN_38[9:0];
    if (sram_even) begin
      if (sizeIsEven) begin
        wmask_0 <= 1'h1;
      end else begin
        if (_T_297) begin
          wmask_0 <= 1'h1;
        end else begin
          if (_T_229) begin
            wmask_0 <= 1'h1;
          end
        end
      end
    end else begin
      if (_T_297) begin
        wmask_0 <= 1'h0;
      end else begin
        if (_T_229) begin
          wmask_0 <= 1'h1;
        end
      end
    end
    if (sram_even) begin
      if (sizeIsEven) begin
        wmask_1 <= 1'h1;
      end else begin
        if (_T_297) begin
          if (_T_299) begin
            wmask_1 <= 1'h0;
          end else begin
            wmask_1 <= 1'h1;
          end
        end else begin
          if (_T_229) begin
            if (_T_356) begin
              wmask_1 <= 1'h0;
            end else begin
              wmask_1 <= 1'h1;
            end
          end
        end
      end
    end else begin
      if (_T_297) begin
        wmask_1 <= 1'h1;
      end else begin
        if (_T_229) begin
          if (_T_439) begin
            wmask_1 <= 1'h0;
          end else begin
            wmask_1 <= 1'h1;
          end
        end
      end
    end
    _T_579 <= io_uop_idx_valid;
    if (_GEN_72) begin
      mem_0_memRead_addr_pipe_0 <= rIdx;
    end
    if (_GEN_72) begin
      mem_1_memRead_addr_pipe_0 <= rIdx;
    end
  end
endmodule
module TensorDataCtrl_2( // @[:@6448.2]
  input          clock, // @[:@6449.4]
  input          io_start, // @[:@6451.4]
  output         io_done, // @[:@6451.4]
  input  [127:0] io_inst, // @[:@6451.4]
  input  [31:0]  io_baddr, // @[:@6451.4]
  input          io_xinit, // @[:@6451.4]
  input          io_xupdate, // @[:@6451.4]
  input          io_yupdate, // @[:@6451.4]
  output         io_stride, // @[:@6451.4]
  output         io_split, // @[:@6451.4]
  output [31:0]  io_addr, // @[:@6451.4]
  output [7:0]   io_len // @[:@6451.4]
);
  wire [31:0] dec_dram_offset; // @[TensorUtil.scala 251:29:@6470.4]
  wire [15:0] dec_ysize; // @[TensorUtil.scala 251:29:@6474.4]
  wire [15:0] dec_xsize; // @[TensorUtil.scala 251:29:@6476.4]
  wire [15:0] dec_xstride; // @[TensorUtil.scala 251:29:@6478.4]
  reg [31:0] caddr; // @[TensorUtil.scala 253:18:@6488.4]
  reg [31:0] _RAND_0;
  reg [31:0] baddr; // @[TensorUtil.scala 254:18:@6489.4]
  reg [31:0] _RAND_1;
  reg [7:0] len; // @[TensorUtil.scala 255:16:@6490.4]
  reg [31:0] _RAND_2;
  reg [7:0] xcnt; // @[TensorUtil.scala 267:17:@6555.4]
  reg [31:0] _RAND_3;
  reg [15:0] xrem; // @[TensorUtil.scala 268:17:@6556.4]
  reg [31:0] _RAND_4;
  wire [18:0] _GEN_27; // @[TensorUtil.scala 269:26:@6557.4]
  wire [18:0] _T_154; // @[TensorUtil.scala 269:26:@6557.4]
  wire [19:0] _T_156; // @[TensorUtil.scala 269:51:@6558.4]
  wire [19:0] _T_157; // @[TensorUtil.scala 269:51:@6559.4]
  wire [18:0] xsize; // @[TensorUtil.scala 269:51:@6560.4]
  reg [15:0] ycnt; // @[TensorUtil.scala 271:17:@6561.4]
  reg [31:0] _RAND_5;
  reg [31:0] xfer_bytes; // @[TensorUtil.scala 273:23:@6562.4]
  reg [31:0] _RAND_6;
  wire [21:0] _GEN_28; // @[TensorUtil.scala 275:35:@6563.4]
  wire [21:0] xstride_bytes; // @[TensorUtil.scala 275:35:@6563.4]
  wire [37:0] _GEN_29; // @[TensorUtil.scala 277:66:@6564.4]
  wire [37:0] _T_160; // @[TensorUtil.scala 277:66:@6564.4]
  wire [37:0] _T_161; // @[TensorUtil.scala 277:47:@6565.4]
  wire [37:0] _GEN_30; // @[TensorUtil.scala 277:33:@6566.4]
  wire [37:0] xfer_init_addr; // @[TensorUtil.scala 277:33:@6566.4]
  wire [32:0] _T_162; // @[TensorUtil.scala 278:31:@6567.4]
  wire [31:0] xfer_split_addr; // @[TensorUtil.scala 278:31:@6568.4]
  wire [31:0] _GEN_31; // @[TensorUtil.scala 279:32:@6569.4]
  wire [32:0] _T_163; // @[TensorUtil.scala 279:32:@6569.4]
  wire [31:0] xfer_stride_addr; // @[TensorUtil.scala 279:32:@6570.4]
  wire [37:0] _GEN_12; // @[TensorUtil.scala 281:55:@6571.4]
  wire [11:0] _T_164; // @[TensorUtil.scala 281:55:@6571.4]
  wire [12:0] _T_165; // @[TensorUtil.scala 281:38:@6572.4]
  wire [12:0] _T_166; // @[TensorUtil.scala 281:38:@6573.4]
  wire [11:0] xfer_init_bytes; // @[TensorUtil.scala 281:38:@6574.4]
  wire [8:0] xfer_init_pulses; // @[TensorUtil.scala 282:43:@6575.4]
  wire [31:0] _GEN_16; // @[TensorUtil.scala 283:56:@6576.4]
  wire [11:0] _T_167; // @[TensorUtil.scala 283:56:@6576.4]
  wire [12:0] _T_168; // @[TensorUtil.scala 283:38:@6577.4]
  wire [12:0] _T_169; // @[TensorUtil.scala 283:38:@6578.4]
  wire [11:0] xfer_split_bytes; // @[TensorUtil.scala 283:38:@6579.4]
  wire [8:0] xfer_split_pulses; // @[TensorUtil.scala 284:44:@6580.4]
  wire [31:0] _GEN_18; // @[TensorUtil.scala 285:57:@6581.4]
  wire [11:0] _T_170; // @[TensorUtil.scala 285:57:@6581.4]
  wire [12:0] _T_171; // @[TensorUtil.scala 285:38:@6582.4]
  wire [12:0] _T_172; // @[TensorUtil.scala 285:38:@6583.4]
  wire [11:0] xfer_stride_bytes; // @[TensorUtil.scala 285:38:@6584.4]
  wire [8:0] xfer_stride_pulses; // @[TensorUtil.scala 286:45:@6585.4]
  wire  _T_173; // @[TensorUtil.scala 288:21:@6586.4]
  wire  _T_175; // @[TensorUtil.scala 289:10:@6587.4]
  wire  _T_176; // @[TensorUtil.scala 288:29:@6588.4]
  wire [16:0] _T_178; // @[TensorUtil.scala 290:24:@6589.4]
  wire [16:0] _T_179; // @[TensorUtil.scala 290:24:@6590.4]
  wire [15:0] _T_180; // @[TensorUtil.scala 290:24:@6591.4]
  wire  _T_181; // @[TensorUtil.scala 290:10:@6592.4]
  wire  stride; // @[TensorUtil.scala 289:18:@6593.4]
  wire  _T_184; // @[TensorUtil.scala 292:35:@6595.4]
  wire  split; // @[TensorUtil.scala 292:28:@6596.4]
  wire [18:0] _GEN_32; // @[TensorUtil.scala 296:16:@6599.6]
  wire  _T_185; // @[TensorUtil.scala 296:16:@6599.6]
  wire [9:0] _T_188; // @[TensorUtil.scala 300:31:@6605.8]
  wire [9:0] _T_189; // @[TensorUtil.scala 300:31:@6606.8]
  wire [8:0] _T_190; // @[TensorUtil.scala 300:31:@6607.8]
  wire [19:0] _T_191; // @[TensorUtil.scala 301:21:@6609.8]
  wire [19:0] _T_192; // @[TensorUtil.scala 301:21:@6610.8]
  wire [18:0] _T_193; // @[TensorUtil.scala 301:21:@6611.8]
  wire [18:0] _GEN_0; // @[TensorUtil.scala 296:36:@6600.6]
  wire [18:0] _GEN_1; // @[TensorUtil.scala 296:36:@6600.6]
  wire  _T_194; // @[TensorUtil.scala 303:25:@6616.6]
  wire [18:0] _GEN_34; // @[TensorUtil.scala 305:16:@6619.8]
  wire  _T_195; // @[TensorUtil.scala 305:16:@6619.8]
  wire [9:0] _T_198; // @[TensorUtil.scala 309:33:@6625.10]
  wire [9:0] _T_199; // @[TensorUtil.scala 309:33:@6626.10]
  wire [8:0] _T_200; // @[TensorUtil.scala 309:33:@6627.10]
  wire [19:0] _T_201; // @[TensorUtil.scala 310:21:@6629.10]
  wire [19:0] _T_202; // @[TensorUtil.scala 310:21:@6630.10]
  wire [18:0] _T_203; // @[TensorUtil.scala 310:21:@6631.10]
  wire [18:0] _GEN_2; // @[TensorUtil.scala 305:38:@6620.8]
  wire [18:0] _GEN_3; // @[TensorUtil.scala 305:38:@6620.8]
  wire  _T_204; // @[TensorUtil.scala 312:25:@6636.8]
  wire [15:0] _GEN_36; // @[TensorUtil.scala 314:15:@6639.10]
  wire  _T_205; // @[TensorUtil.scala 314:15:@6639.10]
  wire [9:0] _T_208; // @[TensorUtil.scala 318:32:@6645.12]
  wire [9:0] _T_209; // @[TensorUtil.scala 318:32:@6646.12]
  wire [8:0] _T_210; // @[TensorUtil.scala 318:32:@6647.12]
  wire [16:0] _T_211; // @[TensorUtil.scala 319:20:@6649.12]
  wire [16:0] _T_212; // @[TensorUtil.scala 319:20:@6650.12]
  wire [15:0] _T_213; // @[TensorUtil.scala 319:20:@6651.12]
  wire [15:0] _GEN_4; // @[TensorUtil.scala 314:36:@6640.10]
  wire [15:0] _GEN_5; // @[TensorUtil.scala 314:36:@6640.10]
  wire [31:0] _GEN_6; // @[TensorUtil.scala 312:35:@6637.8]
  wire [15:0] _GEN_7; // @[TensorUtil.scala 312:35:@6637.8]
  wire [15:0] _GEN_8; // @[TensorUtil.scala 312:35:@6637.8]
  wire [31:0] _GEN_9; // @[TensorUtil.scala 303:36:@6617.6]
  wire [18:0] _GEN_10; // @[TensorUtil.scala 303:36:@6617.6]
  wire [18:0] _GEN_11; // @[TensorUtil.scala 303:36:@6617.6]
  wire [18:0] _GEN_13; // @[TensorUtil.scala 294:18:@6597.4]
  wire [18:0] _GEN_14; // @[TensorUtil.scala 294:18:@6597.4]
  wire [8:0] _T_216; // @[TensorUtil.scala 326:18:@6660.8]
  wire [7:0] _T_217; // @[TensorUtil.scala 326:18:@6661.8]
  wire [7:0] _GEN_15; // @[TensorUtil.scala 325:26:@6659.6]
  wire  _T_219; // @[TensorUtil.scala 331:25:@6668.6]
  wire [16:0] _T_221; // @[TensorUtil.scala 332:18:@6670.8]
  wire [15:0] _T_222; // @[TensorUtil.scala 332:18:@6671.8]
  wire [15:0] _GEN_17; // @[TensorUtil.scala 331:36:@6669.6]
  wire [31:0] _GEN_19; // @[TensorUtil.scala 341:24:@6684.10]
  wire [31:0] _GEN_20; // @[TensorUtil.scala 341:24:@6684.10]
  wire [31:0] _GEN_21; // @[TensorUtil.scala 339:17:@6680.8]
  wire [31:0] _GEN_22; // @[TensorUtil.scala 339:17:@6680.8]
  wire [31:0] _GEN_23; // @[TensorUtil.scala 338:26:@6679.6]
  wire [31:0] _GEN_24; // @[TensorUtil.scala 338:26:@6679.6]
  wire [37:0] _GEN_25; // @[TensorUtil.scala 335:18:@6674.4]
  wire [37:0] _GEN_26; // @[TensorUtil.scala 335:18:@6674.4]
  wire  _T_232; // @[TensorUtil.scala 354:10:@6701.4]
  assign dec_dram_offset = io_inst[56:25]; // @[TensorUtil.scala 251:29:@6470.4]
  assign dec_ysize = io_inst[79:64]; // @[TensorUtil.scala 251:29:@6474.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 251:29:@6476.4]
  assign dec_xstride = io_inst[111:96]; // @[TensorUtil.scala 251:29:@6478.4]
  assign _GEN_27 = {{3'd0}, dec_xsize}; // @[TensorUtil.scala 269:26:@6557.4]
  assign _T_154 = _GEN_27 << 3; // @[TensorUtil.scala 269:26:@6557.4]
  assign _T_156 = _T_154 - 19'h1; // @[TensorUtil.scala 269:51:@6558.4]
  assign _T_157 = $unsigned(_T_156); // @[TensorUtil.scala 269:51:@6559.4]
  assign xsize = _T_157[18:0]; // @[TensorUtil.scala 269:51:@6560.4]
  assign _GEN_28 = {{6'd0}, dec_xstride}; // @[TensorUtil.scala 275:35:@6563.4]
  assign xstride_bytes = _GEN_28 << 6; // @[TensorUtil.scala 275:35:@6563.4]
  assign _GEN_29 = {{6'd0}, dec_dram_offset}; // @[TensorUtil.scala 277:66:@6564.4]
  assign _T_160 = _GEN_29 << 6; // @[TensorUtil.scala 277:66:@6564.4]
  assign _T_161 = 38'hffffffff & _T_160; // @[TensorUtil.scala 277:47:@6565.4]
  assign _GEN_30 = {{6'd0}, io_baddr}; // @[TensorUtil.scala 277:33:@6566.4]
  assign xfer_init_addr = _GEN_30 | _T_161; // @[TensorUtil.scala 277:33:@6566.4]
  assign _T_162 = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@6567.4]
  assign xfer_split_addr = caddr + xfer_bytes; // @[TensorUtil.scala 278:31:@6568.4]
  assign _GEN_31 = {{10'd0}, xstride_bytes}; // @[TensorUtil.scala 279:32:@6569.4]
  assign _T_163 = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@6569.4]
  assign xfer_stride_addr = baddr + _GEN_31; // @[TensorUtil.scala 279:32:@6570.4]
  assign _GEN_12 = xfer_init_addr % 38'h800; // @[TensorUtil.scala 281:55:@6571.4]
  assign _T_164 = _GEN_12[11:0]; // @[TensorUtil.scala 281:55:@6571.4]
  assign _T_165 = 12'h800 - _T_164; // @[TensorUtil.scala 281:38:@6572.4]
  assign _T_166 = $unsigned(_T_165); // @[TensorUtil.scala 281:38:@6573.4]
  assign xfer_init_bytes = _T_166[11:0]; // @[TensorUtil.scala 281:38:@6574.4]
  assign xfer_init_pulses = xfer_init_bytes[11:3]; // @[TensorUtil.scala 282:43:@6575.4]
  assign _GEN_16 = xfer_split_addr % 32'h800; // @[TensorUtil.scala 283:56:@6576.4]
  assign _T_167 = _GEN_16[11:0]; // @[TensorUtil.scala 283:56:@6576.4]
  assign _T_168 = 12'h800 - _T_167; // @[TensorUtil.scala 283:38:@6577.4]
  assign _T_169 = $unsigned(_T_168); // @[TensorUtil.scala 283:38:@6578.4]
  assign xfer_split_bytes = _T_169[11:0]; // @[TensorUtil.scala 283:38:@6579.4]
  assign xfer_split_pulses = xfer_split_bytes[11:3]; // @[TensorUtil.scala 284:44:@6580.4]
  assign _GEN_18 = xfer_stride_addr % 32'h800; // @[TensorUtil.scala 285:57:@6581.4]
  assign _T_170 = _GEN_18[11:0]; // @[TensorUtil.scala 285:57:@6581.4]
  assign _T_171 = 12'h800 - _T_170; // @[TensorUtil.scala 285:38:@6582.4]
  assign _T_172 = $unsigned(_T_171); // @[TensorUtil.scala 285:38:@6583.4]
  assign xfer_stride_bytes = _T_172[11:0]; // @[TensorUtil.scala 285:38:@6584.4]
  assign xfer_stride_pulses = xfer_stride_bytes[11:3]; // @[TensorUtil.scala 286:45:@6585.4]
  assign _T_173 = xcnt == len; // @[TensorUtil.scala 288:21:@6586.4]
  assign _T_175 = xrem == 16'h0; // @[TensorUtil.scala 289:10:@6587.4]
  assign _T_176 = _T_173 & _T_175; // @[TensorUtil.scala 288:29:@6588.4]
  assign _T_178 = dec_ysize - 16'h1; // @[TensorUtil.scala 290:24:@6589.4]
  assign _T_179 = $unsigned(_T_178); // @[TensorUtil.scala 290:24:@6590.4]
  assign _T_180 = _T_179[15:0]; // @[TensorUtil.scala 290:24:@6591.4]
  assign _T_181 = ycnt != _T_180; // @[TensorUtil.scala 290:10:@6592.4]
  assign stride = _T_176 & _T_181; // @[TensorUtil.scala 289:18:@6593.4]
  assign _T_184 = xrem != 16'h0; // @[TensorUtil.scala 292:35:@6595.4]
  assign split = _T_173 & _T_184; // @[TensorUtil.scala 292:28:@6596.4]
  assign _GEN_32 = {{10'd0}, xfer_init_pulses}; // @[TensorUtil.scala 296:16:@6599.6]
  assign _T_185 = xsize < _GEN_32; // @[TensorUtil.scala 296:16:@6599.6]
  assign _T_188 = xfer_init_pulses - 9'h1; // @[TensorUtil.scala 300:31:@6605.8]
  assign _T_189 = $unsigned(_T_188); // @[TensorUtil.scala 300:31:@6606.8]
  assign _T_190 = _T_189[8:0]; // @[TensorUtil.scala 300:31:@6607.8]
  assign _T_191 = xsize - _GEN_32; // @[TensorUtil.scala 301:21:@6609.8]
  assign _T_192 = $unsigned(_T_191); // @[TensorUtil.scala 301:21:@6610.8]
  assign _T_193 = _T_192[18:0]; // @[TensorUtil.scala 301:21:@6611.8]
  assign _GEN_0 = _T_185 ? xsize : {{10'd0}, _T_190}; // @[TensorUtil.scala 296:36:@6600.6]
  assign _GEN_1 = _T_185 ? 19'h0 : _T_193; // @[TensorUtil.scala 296:36:@6600.6]
  assign _T_194 = io_xupdate & stride; // @[TensorUtil.scala 303:25:@6616.6]
  assign _GEN_34 = {{10'd0}, xfer_stride_pulses}; // @[TensorUtil.scala 305:16:@6619.8]
  assign _T_195 = xsize < _GEN_34; // @[TensorUtil.scala 305:16:@6619.8]
  assign _T_198 = xfer_stride_pulses - 9'h1; // @[TensorUtil.scala 309:33:@6625.10]
  assign _T_199 = $unsigned(_T_198); // @[TensorUtil.scala 309:33:@6626.10]
  assign _T_200 = _T_199[8:0]; // @[TensorUtil.scala 309:33:@6627.10]
  assign _T_201 = xsize - _GEN_34; // @[TensorUtil.scala 310:21:@6629.10]
  assign _T_202 = $unsigned(_T_201); // @[TensorUtil.scala 310:21:@6630.10]
  assign _T_203 = _T_202[18:0]; // @[TensorUtil.scala 310:21:@6631.10]
  assign _GEN_2 = _T_195 ? xsize : {{10'd0}, _T_200}; // @[TensorUtil.scala 305:38:@6620.8]
  assign _GEN_3 = _T_195 ? 19'h0 : _T_203; // @[TensorUtil.scala 305:38:@6620.8]
  assign _T_204 = io_xupdate & split; // @[TensorUtil.scala 312:25:@6636.8]
  assign _GEN_36 = {{7'd0}, xfer_split_pulses}; // @[TensorUtil.scala 314:15:@6639.10]
  assign _T_205 = xrem < _GEN_36; // @[TensorUtil.scala 314:15:@6639.10]
  assign _T_208 = xfer_split_pulses - 9'h1; // @[TensorUtil.scala 318:32:@6645.12]
  assign _T_209 = $unsigned(_T_208); // @[TensorUtil.scala 318:32:@6646.12]
  assign _T_210 = _T_209[8:0]; // @[TensorUtil.scala 318:32:@6647.12]
  assign _T_211 = xrem - _GEN_36; // @[TensorUtil.scala 319:20:@6649.12]
  assign _T_212 = $unsigned(_T_211); // @[TensorUtil.scala 319:20:@6650.12]
  assign _T_213 = _T_212[15:0]; // @[TensorUtil.scala 319:20:@6651.12]
  assign _GEN_4 = _T_205 ? xrem : {{7'd0}, _T_210}; // @[TensorUtil.scala 314:36:@6640.10]
  assign _GEN_5 = _T_205 ? 16'h0 : _T_213; // @[TensorUtil.scala 314:36:@6640.10]
  assign _GEN_6 = _T_204 ? {{20'd0}, xfer_split_bytes} : xfer_bytes; // @[TensorUtil.scala 312:35:@6637.8]
  assign _GEN_7 = _T_204 ? _GEN_4 : {{8'd0}, len}; // @[TensorUtil.scala 312:35:@6637.8]
  assign _GEN_8 = _T_204 ? _GEN_5 : xrem; // @[TensorUtil.scala 312:35:@6637.8]
  assign _GEN_9 = _T_194 ? {{20'd0}, xfer_stride_bytes} : _GEN_6; // @[TensorUtil.scala 303:36:@6617.6]
  assign _GEN_10 = _T_194 ? _GEN_2 : {{3'd0}, _GEN_7}; // @[TensorUtil.scala 303:36:@6617.6]
  assign _GEN_11 = _T_194 ? _GEN_3 : {{3'd0}, _GEN_8}; // @[TensorUtil.scala 303:36:@6617.6]
  assign _GEN_13 = io_start ? _GEN_0 : _GEN_10; // @[TensorUtil.scala 294:18:@6597.4]
  assign _GEN_14 = io_start ? _GEN_1 : _GEN_11; // @[TensorUtil.scala 294:18:@6597.4]
  assign _T_216 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@6660.8]
  assign _T_217 = xcnt + 8'h1; // @[TensorUtil.scala 326:18:@6661.8]
  assign _GEN_15 = io_xupdate ? _T_217 : xcnt; // @[TensorUtil.scala 325:26:@6659.6]
  assign _T_219 = io_yupdate & stride; // @[TensorUtil.scala 331:25:@6668.6]
  assign _T_221 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@6670.8]
  assign _T_222 = ycnt + 16'h1; // @[TensorUtil.scala 332:18:@6671.8]
  assign _GEN_17 = _T_219 ? _T_222 : ycnt; // @[TensorUtil.scala 331:36:@6669.6]
  assign _GEN_19 = stride ? xfer_stride_addr : caddr; // @[TensorUtil.scala 341:24:@6684.10]
  assign _GEN_20 = stride ? xfer_stride_addr : baddr; // @[TensorUtil.scala 341:24:@6684.10]
  assign _GEN_21 = split ? xfer_split_addr : _GEN_19; // @[TensorUtil.scala 339:17:@6680.8]
  assign _GEN_22 = split ? baddr : _GEN_20; // @[TensorUtil.scala 339:17:@6680.8]
  assign _GEN_23 = io_yupdate ? _GEN_21 : caddr; // @[TensorUtil.scala 338:26:@6679.6]
  assign _GEN_24 = io_yupdate ? _GEN_22 : baddr; // @[TensorUtil.scala 338:26:@6679.6]
  assign _GEN_25 = io_start ? xfer_init_addr : {{6'd0}, _GEN_23}; // @[TensorUtil.scala 335:18:@6674.4]
  assign _GEN_26 = io_start ? xfer_init_addr : {{6'd0}, _GEN_24}; // @[TensorUtil.scala 335:18:@6674.4]
  assign _T_232 = ycnt == _T_180; // @[TensorUtil.scala 354:10:@6701.4]
  assign io_done = _T_176 & _T_232; // @[TensorUtil.scala 352:11:@6703.4]
  assign io_stride = _T_176 & _T_181; // @[TensorUtil.scala 347:13:@6689.4]
  assign io_split = _T_173 & _T_184; // @[TensorUtil.scala 348:12:@6690.4]
  assign io_addr = caddr; // @[TensorUtil.scala 350:11:@6693.4]
  assign io_len = len; // @[TensorUtil.scala 351:10:@6694.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  caddr = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  baddr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  len = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  xcnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xrem = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ycnt = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  xfer_bytes = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    caddr <= _GEN_25[31:0];
    baddr <= _GEN_26[31:0];
    len <= _GEN_13[7:0];
    if (io_xinit) begin
      xcnt <= 8'h0;
    end else begin
      if (io_xupdate) begin
        xcnt <= _T_217;
      end
    end
    xrem <= _GEN_14[15:0];
    if (io_start) begin
      ycnt <= 16'h0;
    end else begin
      if (_T_219) begin
        ycnt <= _T_222;
      end
    end
    if (io_start) begin
      xfer_bytes <= {{20'd0}, xfer_init_bytes};
    end else begin
      if (_T_194) begin
        xfer_bytes <= {{20'd0}, xfer_stride_bytes};
      end else begin
        if (_T_204) begin
          xfer_bytes <= {{20'd0}, xfer_split_bytes};
        end
      end
    end
  end
endmodule
module TensorPadCtrl_8( // @[:@6705.2]
  input          clock, // @[:@6706.4]
  input          reset, // @[:@6707.4]
  input          io_start, // @[:@6708.4]
  output         io_done, // @[:@6708.4]
  input  [127:0] io_inst // @[:@6708.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@6733.4]
  wire [3:0] dec_ypad_0; // @[TensorUtil.scala 173:29:@6737.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@6741.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@6743.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@6745.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@6746.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@6747.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@6748.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@6749.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@6749.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@6750.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@6751.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@6751.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@6752.4]
  wire [18:0] _GEN_12; // @[TensorUtil.scala 182:46:@6753.4]
  wire [18:0] _T_39; // @[TensorUtil.scala 182:46:@6753.4]
  wire [19:0] _T_41; // @[TensorUtil.scala 182:71:@6754.4]
  wire [19:0] _T_42; // @[TensorUtil.scala 182:71:@6755.4]
  wire [18:0] xval; // @[TensorUtil.scala 182:71:@6756.4]
  wire  _T_44; // @[TensorUtil.scala 190:22:@6757.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 190:42:@6758.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 190:42:@6759.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 190:42:@6760.4]
  wire [3:0] yval; // @[TensorUtil.scala 190:10:@6761.4]
  reg  state; // @[TensorUtil.scala 197:22:@6762.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@6763.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@6765.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@6772.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@6773.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@6774.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@6775.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@6771.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@6764.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@6779.4]
  wire [18:0] _GEN_4; // @[TensorUtil.scala 212:25:@6780.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@6786.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@6793.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@6794.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@6792.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@6798.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@6799.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@6806.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@6808.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@6809.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@6807.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@6814.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@6733.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorUtil.scala 173:29:@6737.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@6741.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@6743.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@6749.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@6749.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@6750.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@6751.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@6751.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@6752.4]
  assign _GEN_12 = {{3'd0}, _T_38}; // @[TensorUtil.scala 182:46:@6753.4]
  assign _T_39 = _GEN_12 << 3; // @[TensorUtil.scala 182:46:@6753.4]
  assign _T_41 = _T_39 - 19'h1; // @[TensorUtil.scala 182:71:@6754.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@6755.4]
  assign xval = _T_42[18:0]; // @[TensorUtil.scala 182:71:@6756.4]
  assign _T_44 = dec_ypad_0 != 4'h0; // @[TensorUtil.scala 190:22:@6757.4]
  assign _T_46 = dec_ypad_0 - 4'h1; // @[TensorUtil.scala 190:42:@6758.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 190:42:@6759.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 190:42:@6760.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 190:10:@6761.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@6763.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@6765.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@6772.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@6773.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@6774.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@6775.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@6771.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@6764.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@6779.4]
  assign _GEN_4 = _T_56 ? xval : {{3'd0}, xmax}; // @[TensorUtil.scala 212:25:@6780.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@6786.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6793.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6794.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@6792.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@6798.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@6799.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@6806.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@6808.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@6809.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@6807.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@6814.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@6817.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_9( // @[:@6819.2]
  input          clock, // @[:@6820.4]
  input          reset, // @[:@6821.4]
  input          io_start, // @[:@6822.4]
  output         io_done, // @[:@6822.4]
  input  [127:0] io_inst // @[:@6822.4]
);
  wire [15:0] dec_xsize; // @[TensorUtil.scala 173:29:@6847.4]
  wire [3:0] dec_ypad_1; // @[TensorUtil.scala 173:29:@6853.4]
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@6855.4]
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@6857.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@6859.4]
  reg [31:0] _RAND_0;
  reg [3:0] ymax; // @[TensorUtil.scala 176:17:@6860.4]
  reg [31:0] _RAND_1;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@6861.4]
  reg [31:0] _RAND_2;
  reg [3:0] ycnt; // @[TensorUtil.scala 178:17:@6862.4]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_10; // @[TensorUtil.scala 182:20:@6863.4]
  wire [16:0] _T_35; // @[TensorUtil.scala 182:20:@6863.4]
  wire [15:0] _T_36; // @[TensorUtil.scala 182:20:@6864.4]
  wire [15:0] _GEN_11; // @[TensorUtil.scala 182:32:@6865.4]
  wire [16:0] _T_37; // @[TensorUtil.scala 182:32:@6865.4]
  wire [15:0] _T_38; // @[TensorUtil.scala 182:32:@6866.4]
  wire [18:0] _GEN_12; // @[TensorUtil.scala 182:46:@6867.4]
  wire [18:0] _T_39; // @[TensorUtil.scala 182:46:@6867.4]
  wire [19:0] _T_41; // @[TensorUtil.scala 182:71:@6868.4]
  wire [19:0] _T_42; // @[TensorUtil.scala 182:71:@6869.4]
  wire [18:0] xval; // @[TensorUtil.scala 182:71:@6870.4]
  wire  _T_44; // @[TensorUtil.scala 192:22:@6871.4]
  wire [4:0] _T_46; // @[TensorUtil.scala 192:42:@6872.4]
  wire [4:0] _T_47; // @[TensorUtil.scala 192:42:@6873.4]
  wire [3:0] _T_48; // @[TensorUtil.scala 192:42:@6874.4]
  wire [3:0] yval; // @[TensorUtil.scala 192:10:@6875.4]
  reg  state; // @[TensorUtil.scala 197:22:@6876.4]
  reg [31:0] _RAND_4;
  wire  _T_51; // @[Conditional.scala 37:30:@6877.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@6879.6]
  wire  _T_53; // @[TensorUtil.scala 206:17:@6886.8]
  wire  _T_54; // @[TensorUtil.scala 206:34:@6887.8]
  wire  _T_55; // @[TensorUtil.scala 206:26:@6888.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@6889.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@6885.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@6878.4]
  wire  _T_56; // @[TensorUtil.scala 212:14:@6893.4]
  wire [18:0] _GEN_4; // @[TensorUtil.scala 212:25:@6894.4]
  wire  _T_59; // @[TensorUtil.scala 217:24:@6900.4]
  wire [16:0] _T_63; // @[TensorUtil.scala 220:18:@6907.8]
  wire [15:0] _T_64; // @[TensorUtil.scala 220:18:@6908.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@6906.6]
  wire  _T_67; // @[TensorUtil.scala 223:32:@6912.4]
  wire  _T_68; // @[TensorUtil.scala 223:24:@6913.4]
  wire  _T_72; // @[TensorUtil.scala 225:32:@6920.6]
  wire [4:0] _T_74; // @[TensorUtil.scala 226:18:@6922.8]
  wire [3:0] _T_75; // @[TensorUtil.scala 226:18:@6923.8]
  wire [3:0] _GEN_8; // @[TensorUtil.scala 225:50:@6921.6]
  wire  _T_78; // @[TensorUtil.scala 229:32:@6928.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorUtil.scala 173:29:@6847.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorUtil.scala 173:29:@6853.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@6855.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@6857.4]
  assign _GEN_10 = {{12'd0}, dec_xpad_0}; // @[TensorUtil.scala 182:20:@6863.4]
  assign _T_35 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@6863.4]
  assign _T_36 = _GEN_10 + dec_xsize; // @[TensorUtil.scala 182:20:@6864.4]
  assign _GEN_11 = {{12'd0}, dec_xpad_1}; // @[TensorUtil.scala 182:32:@6865.4]
  assign _T_37 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@6865.4]
  assign _T_38 = _T_36 + _GEN_11; // @[TensorUtil.scala 182:32:@6866.4]
  assign _GEN_12 = {{3'd0}, _T_38}; // @[TensorUtil.scala 182:46:@6867.4]
  assign _T_39 = _GEN_12 << 3; // @[TensorUtil.scala 182:46:@6867.4]
  assign _T_41 = _T_39 - 19'h1; // @[TensorUtil.scala 182:71:@6868.4]
  assign _T_42 = $unsigned(_T_41); // @[TensorUtil.scala 182:71:@6869.4]
  assign xval = _T_42[18:0]; // @[TensorUtil.scala 182:71:@6870.4]
  assign _T_44 = dec_ypad_1 != 4'h0; // @[TensorUtil.scala 192:22:@6871.4]
  assign _T_46 = dec_ypad_1 - 4'h1; // @[TensorUtil.scala 192:42:@6872.4]
  assign _T_47 = $unsigned(_T_46); // @[TensorUtil.scala 192:42:@6873.4]
  assign _T_48 = _T_47[3:0]; // @[TensorUtil.scala 192:42:@6874.4]
  assign yval = _T_44 ? _T_48 : 4'h0; // @[TensorUtil.scala 192:10:@6875.4]
  assign _T_51 = 1'h0 == state; // @[Conditional.scala 37:30:@6877.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@6879.6]
  assign _T_53 = ycnt == ymax; // @[TensorUtil.scala 206:17:@6886.8]
  assign _T_54 = xcnt == xmax; // @[TensorUtil.scala 206:34:@6887.8]
  assign _T_55 = _T_53 & _T_54; // @[TensorUtil.scala 206:26:@6888.8]
  assign _GEN_1 = _T_55 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@6889.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@6885.6]
  assign _GEN_3 = _T_51 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@6878.4]
  assign _T_56 = state == 1'h0; // @[TensorUtil.scala 212:14:@6893.4]
  assign _GEN_4 = _T_56 ? xval : {{3'd0}, xmax}; // @[TensorUtil.scala 212:25:@6894.4]
  assign _T_59 = _T_56 | _T_54; // @[TensorUtil.scala 217:24:@6900.4]
  assign _T_63 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6907.8]
  assign _T_64 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@6908.8]
  assign _GEN_6 = state ? _T_64 : xcnt; // @[TensorUtil.scala 219:33:@6906.6]
  assign _T_67 = ymax == 4'h0; // @[TensorUtil.scala 223:32:@6912.4]
  assign _T_68 = _T_56 | _T_67; // @[TensorUtil.scala 223:24:@6913.4]
  assign _T_72 = state & _T_54; // @[TensorUtil.scala 225:32:@6920.6]
  assign _T_74 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@6922.8]
  assign _T_75 = ycnt + 4'h1; // @[TensorUtil.scala 226:18:@6923.8]
  assign _GEN_8 = _T_72 ? _T_75 : ycnt; // @[TensorUtil.scala 225:50:@6921.6]
  assign _T_78 = state & _T_53; // @[TensorUtil.scala 229:32:@6928.4]
  assign io_done = _T_78 & _T_54; // @[TensorUtil.scala 229:11:@6931.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ymax = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  xcnt = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ycnt = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    xmax <= _GEN_4[15:0];
    if (_T_56) begin
      if (_T_44) begin
        ymax <= _T_48;
      end else begin
        ymax <= 4'h0;
      end
    end
    if (_T_59) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_64;
      end
    end
    if (_T_68) begin
      ycnt <= 4'h0;
    end else begin
      if (_T_72) begin
        ycnt <= _T_75;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_51) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_10( // @[:@6933.2]
  input          clock, // @[:@6934.4]
  input          reset, // @[:@6935.4]
  input          io_start, // @[:@6936.4]
  output         io_done, // @[:@6936.4]
  input  [127:0] io_inst // @[:@6936.4]
);
  wire [3:0] dec_xpad_0; // @[TensorUtil.scala 173:29:@6969.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@6973.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@6975.4]
  reg [31:0] _RAND_1;
  wire [6:0] _GEN_10; // @[TensorUtil.scala 184:19:@6977.4]
  wire [6:0] _T_35; // @[TensorUtil.scala 184:19:@6977.4]
  wire [7:0] _T_37; // @[TensorUtil.scala 184:44:@6978.4]
  wire [7:0] _T_38; // @[TensorUtil.scala 184:44:@6979.4]
  wire [6:0] xval; // @[TensorUtil.scala 184:44:@6980.4]
  reg  state; // @[TensorUtil.scala 197:22:@6981.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@6982.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@6984.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@6992.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@6994.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@6990.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@6983.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@6998.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@7005.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@7012.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@7013.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@7011.6]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorUtil.scala 173:29:@6969.4]
  assign _GEN_10 = {{3'd0}, dec_xpad_0}; // @[TensorUtil.scala 184:19:@6977.4]
  assign _T_35 = _GEN_10 << 3; // @[TensorUtil.scala 184:19:@6977.4]
  assign _T_37 = _T_35 - 7'h1; // @[TensorUtil.scala 184:44:@6978.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 184:44:@6979.4]
  assign xval = _T_38[6:0]; // @[TensorUtil.scala 184:44:@6980.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@6982.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@6984.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@6992.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@6994.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@6990.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@6983.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@6998.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@7005.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@7012.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@7013.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@7011.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@7036.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{9'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorPadCtrl_11( // @[:@7038.2]
  input          clock, // @[:@7039.4]
  input          reset, // @[:@7040.4]
  input          io_start, // @[:@7041.4]
  output         io_done, // @[:@7041.4]
  input  [127:0] io_inst // @[:@7041.4]
);
  wire [3:0] dec_xpad_1; // @[TensorUtil.scala 173:29:@7076.4]
  reg [15:0] xmax; // @[TensorUtil.scala 175:17:@7078.4]
  reg [31:0] _RAND_0;
  reg [15:0] xcnt; // @[TensorUtil.scala 177:17:@7080.4]
  reg [31:0] _RAND_1;
  wire [6:0] _GEN_10; // @[TensorUtil.scala 186:19:@7082.4]
  wire [6:0] _T_35; // @[TensorUtil.scala 186:19:@7082.4]
  wire [7:0] _T_37; // @[TensorUtil.scala 186:44:@7083.4]
  wire [7:0] _T_38; // @[TensorUtil.scala 186:44:@7084.4]
  wire [6:0] xval; // @[TensorUtil.scala 186:44:@7085.4]
  reg  state; // @[TensorUtil.scala 197:22:@7086.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[Conditional.scala 37:30:@7087.4]
  wire  _GEN_0; // @[TensorUtil.scala 201:22:@7089.6]
  wire  _T_43; // @[TensorUtil.scala 206:34:@7097.8]
  wire  _GEN_1; // @[TensorUtil.scala 206:44:@7099.8]
  wire  _GEN_2; // @[Conditional.scala 39:67:@7095.6]
  wire  _GEN_3; // @[Conditional.scala 40:58:@7088.4]
  wire  _T_45; // @[TensorUtil.scala 212:14:@7103.4]
  wire  _T_48; // @[TensorUtil.scala 217:24:@7110.4]
  wire [16:0] _T_52; // @[TensorUtil.scala 220:18:@7117.8]
  wire [15:0] _T_53; // @[TensorUtil.scala 220:18:@7118.8]
  wire [15:0] _GEN_6; // @[TensorUtil.scala 219:33:@7116.6]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorUtil.scala 173:29:@7076.4]
  assign _GEN_10 = {{3'd0}, dec_xpad_1}; // @[TensorUtil.scala 186:19:@7082.4]
  assign _T_35 = _GEN_10 << 3; // @[TensorUtil.scala 186:19:@7082.4]
  assign _T_37 = _T_35 - 7'h1; // @[TensorUtil.scala 186:44:@7083.4]
  assign _T_38 = $unsigned(_T_37); // @[TensorUtil.scala 186:44:@7084.4]
  assign xval = _T_38[6:0]; // @[TensorUtil.scala 186:44:@7085.4]
  assign _T_40 = 1'h0 == state; // @[Conditional.scala 37:30:@7087.4]
  assign _GEN_0 = io_start ? 1'h1 : state; // @[TensorUtil.scala 201:22:@7089.6]
  assign _T_43 = xcnt == xmax; // @[TensorUtil.scala 206:34:@7097.8]
  assign _GEN_1 = _T_43 ? 1'h0 : state; // @[TensorUtil.scala 206:44:@7099.8]
  assign _GEN_2 = state ? _GEN_1 : state; // @[Conditional.scala 39:67:@7095.6]
  assign _GEN_3 = _T_40 ? _GEN_0 : _GEN_2; // @[Conditional.scala 40:58:@7088.4]
  assign _T_45 = state == 1'h0; // @[TensorUtil.scala 212:14:@7103.4]
  assign _T_48 = _T_45 | _T_43; // @[TensorUtil.scala 217:24:@7110.4]
  assign _T_52 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@7117.8]
  assign _T_53 = xcnt + 16'h1; // @[TensorUtil.scala 220:18:@7118.8]
  assign _GEN_6 = state ? _T_53 : xcnt; // @[TensorUtil.scala 219:33:@7116.6]
  assign io_done = state & _T_43; // @[TensorUtil.scala 229:11:@7141.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  xmax = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  xcnt = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_45) begin
      xmax <= {{9'd0}, xval};
    end
    if (_T_48) begin
      xcnt <= 16'h0;
    end else begin
      if (state) begin
        xcnt <= _T_53;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_40) begin
        if (io_start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_43) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module TensorLoad_2( // @[:@7143.2]
  input          clock, // @[:@7144.4]
  input          reset, // @[:@7145.4]
  input          io_start, // @[:@7146.4]
  output         io_done, // @[:@7146.4]
  input  [127:0] io_inst, // @[:@7146.4]
  input  [31:0]  io_baddr, // @[:@7146.4]
  input          io_vme_rd_cmd_ready, // @[:@7146.4]
  output         io_vme_rd_cmd_valid, // @[:@7146.4]
  output [31:0]  io_vme_rd_cmd_bits_addr, // @[:@7146.4]
  output [7:0]   io_vme_rd_cmd_bits_len, // @[:@7146.4]
  output         io_vme_rd_data_ready, // @[:@7146.4]
  input          io_vme_rd_data_valid, // @[:@7146.4]
  input  [63:0]  io_vme_rd_data_bits, // @[:@7146.4]
  input          io_tensor_rd_idx_valid, // @[:@7146.4]
  input  [10:0]  io_tensor_rd_idx_bits, // @[:@7146.4]
  output         io_tensor_rd_data_valid, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_0, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_1, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_2, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_3, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_4, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_5, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_6, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_7, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_8, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_9, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_10, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_11, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_12, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_13, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_14, // @[:@7146.4]
  output [31:0]  io_tensor_rd_data_bits_0_15, // @[:@7146.4]
  input          io_tensor_wr_valid, // @[:@7146.4]
  input  [10:0]  io_tensor_wr_bits_idx, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_0, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_1, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_2, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_3, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_4, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_5, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_6, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_7, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_8, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_9, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_10, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_11, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_12, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_13, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_14, // @[:@7146.4]
  input  [31:0]  io_tensor_wr_bits_data_0_15 // @[:@7146.4]
);
  wire  dataCtrl_clock; // @[TensorLoad.scala 52:24:@7183.4]
  wire  dataCtrl_io_start; // @[TensorLoad.scala 52:24:@7183.4]
  wire  dataCtrl_io_done; // @[TensorLoad.scala 52:24:@7183.4]
  wire [127:0] dataCtrl_io_inst; // @[TensorLoad.scala 52:24:@7183.4]
  wire [31:0] dataCtrl_io_baddr; // @[TensorLoad.scala 52:24:@7183.4]
  wire  dataCtrl_io_xinit; // @[TensorLoad.scala 52:24:@7183.4]
  wire  dataCtrl_io_xupdate; // @[TensorLoad.scala 52:24:@7183.4]
  wire  dataCtrl_io_yupdate; // @[TensorLoad.scala 52:24:@7183.4]
  wire  dataCtrl_io_stride; // @[TensorLoad.scala 52:24:@7183.4]
  wire  dataCtrl_io_split; // @[TensorLoad.scala 52:24:@7183.4]
  wire [31:0] dataCtrl_io_addr; // @[TensorLoad.scala 52:24:@7183.4]
  wire [7:0] dataCtrl_io_len; // @[TensorLoad.scala 52:24:@7183.4]
  wire  yPadCtrl0_clock; // @[TensorLoad.scala 55:25:@7187.4]
  wire  yPadCtrl0_reset; // @[TensorLoad.scala 55:25:@7187.4]
  wire  yPadCtrl0_io_start; // @[TensorLoad.scala 55:25:@7187.4]
  wire  yPadCtrl0_io_done; // @[TensorLoad.scala 55:25:@7187.4]
  wire [127:0] yPadCtrl0_io_inst; // @[TensorLoad.scala 55:25:@7187.4]
  wire  yPadCtrl1_clock; // @[TensorLoad.scala 56:25:@7190.4]
  wire  yPadCtrl1_reset; // @[TensorLoad.scala 56:25:@7190.4]
  wire  yPadCtrl1_io_start; // @[TensorLoad.scala 56:25:@7190.4]
  wire  yPadCtrl1_io_done; // @[TensorLoad.scala 56:25:@7190.4]
  wire [127:0] yPadCtrl1_io_inst; // @[TensorLoad.scala 56:25:@7190.4]
  wire  xPadCtrl0_clock; // @[TensorLoad.scala 57:25:@7193.4]
  wire  xPadCtrl0_reset; // @[TensorLoad.scala 57:25:@7193.4]
  wire  xPadCtrl0_io_start; // @[TensorLoad.scala 57:25:@7193.4]
  wire  xPadCtrl0_io_done; // @[TensorLoad.scala 57:25:@7193.4]
  wire [127:0] xPadCtrl0_io_inst; // @[TensorLoad.scala 57:25:@7193.4]
  wire  xPadCtrl1_clock; // @[TensorLoad.scala 58:25:@7196.4]
  wire  xPadCtrl1_reset; // @[TensorLoad.scala 58:25:@7196.4]
  wire  xPadCtrl1_io_start; // @[TensorLoad.scala 58:25:@7196.4]
  wire  xPadCtrl1_io_done; // @[TensorLoad.scala 58:25:@7196.4]
  wire [127:0] xPadCtrl1_io_inst; // @[TensorLoad.scala 58:25:@7196.4]
  reg [63:0] tensorFile_0_0 [0:2047]; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] _RAND_0;
  wire [63:0] tensorFile_0_0_rdata_0_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_0_rdata_0_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire [63:0] tensorFile_0_0__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_0__T_992_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_0__T_992_mask; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_0__T_992_en; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] tensorFile_0_1 [0:2047]; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] _RAND_1;
  wire [63:0] tensorFile_0_1_rdata_0_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_1_rdata_0_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire [63:0] tensorFile_0_1__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_1__T_992_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_1__T_992_mask; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_1__T_992_en; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] tensorFile_0_2 [0:2047]; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] _RAND_2;
  wire [63:0] tensorFile_0_2_rdata_0_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_2_rdata_0_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire [63:0] tensorFile_0_2__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_2__T_992_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_2__T_992_mask; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_2__T_992_en; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] tensorFile_0_3 [0:2047]; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] _RAND_3;
  wire [63:0] tensorFile_0_3_rdata_0_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_3_rdata_0_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire [63:0] tensorFile_0_3__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_3__T_992_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_3__T_992_mask; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_3__T_992_en; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] tensorFile_0_4 [0:2047]; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] _RAND_4;
  wire [63:0] tensorFile_0_4_rdata_0_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_4_rdata_0_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire [63:0] tensorFile_0_4__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_4__T_992_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_4__T_992_mask; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_4__T_992_en; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] tensorFile_0_5 [0:2047]; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] _RAND_5;
  wire [63:0] tensorFile_0_5_rdata_0_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_5_rdata_0_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire [63:0] tensorFile_0_5__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_5__T_992_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_5__T_992_mask; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_5__T_992_en; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] tensorFile_0_6 [0:2047]; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] _RAND_6;
  wire [63:0] tensorFile_0_6_rdata_0_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_6_rdata_0_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire [63:0] tensorFile_0_6__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_6__T_992_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_6__T_992_mask; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_6__T_992_en; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] tensorFile_0_7 [0:2047]; // @[TensorLoad.scala 222:16:@7466.4]
  reg [63:0] _RAND_7;
  wire [63:0] tensorFile_0_7_rdata_0_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_7_rdata_0_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire [63:0] tensorFile_0_7__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
  wire [10:0] tensorFile_0_7__T_992_addr; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_7__T_992_mask; // @[TensorLoad.scala 222:16:@7466.4]
  wire  tensorFile_0_7__T_992_en; // @[TensorLoad.scala 222:16:@7466.4]
  wire [15:0] dec_sram_offset; // @[TensorLoad.scala 51:29:@7163.4]
  wire [15:0] dec_xsize; // @[TensorLoad.scala 51:29:@7171.4]
  wire [3:0] dec_ypad_0; // @[TensorLoad.scala 51:29:@7175.4]
  wire [3:0] dec_ypad_1; // @[TensorLoad.scala 51:29:@7177.4]
  wire [3:0] dec_xpad_0; // @[TensorLoad.scala 51:29:@7179.4]
  wire [3:0] dec_xpad_1; // @[TensorLoad.scala 51:29:@7181.4]
  reg  dataCtrlDone; // @[TensorLoad.scala 54:29:@7186.4]
  reg [31:0] _RAND_8;
  reg [2:0] tag; // @[TensorLoad.scala 60:16:@7199.4]
  reg [31:0] _RAND_9;
  reg [2:0] state; // @[TensorLoad.scala 65:22:@7201.4]
  reg [31:0] _RAND_10;
  wire  _T_614; // @[Conditional.scala 37:30:@7202.4]
  wire  _T_616; // @[TensorLoad.scala 71:25:@7205.8]
  wire  _T_618; // @[TensorLoad.scala 73:31:@7210.10]
  wire [2:0] _GEN_0; // @[TensorLoad.scala 73:40:@7211.10]
  wire [2:0] _GEN_1; // @[TensorLoad.scala 71:34:@7206.8]
  wire [2:0] _GEN_2; // @[TensorLoad.scala 70:22:@7204.6]
  wire  _T_619; // @[Conditional.scala 37:30:@7220.6]
  wire [2:0] _GEN_4; // @[TensorLoad.scala 81:31:@7222.8]
  wire  _T_622; // @[Conditional.scala 37:30:@7233.8]
  wire [2:0] _GEN_5; // @[TensorLoad.scala 90:31:@7235.10]
  wire  _T_623; // @[Conditional.scala 37:30:@7240.10]
  wire [2:0] _GEN_6; // @[TensorLoad.scala 95:33:@7242.12]
  wire  _T_624; // @[Conditional.scala 37:30:@7247.12]
  wire  _T_626; // @[TensorLoad.scala 102:27:@7251.18]
  wire  _T_628; // @[TensorLoad.scala 104:33:@7256.20]
  wire [2:0] _GEN_7; // @[TensorLoad.scala 104:42:@7257.20]
  wire [2:0] _GEN_8; // @[TensorLoad.scala 102:36:@7252.18]
  wire [2:0] _GEN_10; // @[TensorLoad.scala 110:36:@7267.20]
  wire [2:0] _GEN_11; // @[TensorLoad.scala 117:39:@7280.20]
  wire [2:0] _GEN_12; // @[TensorLoad.scala 109:40:@7265.18]
  wire [2:0] _GEN_13; // @[TensorLoad.scala 101:32:@7250.16]
  wire [2:0] _GEN_14; // @[TensorLoad.scala 100:34:@7249.14]
  wire  _T_633; // @[Conditional.scala 37:30:@7286.14]
  wire [2:0] _GEN_17; // @[TensorLoad.scala 124:28:@7289.18]
  wire [2:0] _GEN_18; // @[TensorLoad.scala 123:31:@7288.16]
  wire  _T_638; // @[Conditional.scala 37:30:@7310.16]
  wire  _T_639; // @[TensorLoad.scala 140:30:@7312.18]
  wire [2:0] _GEN_19; // @[TensorLoad.scala 140:47:@7313.18]
  wire [2:0] _GEN_20; // @[Conditional.scala 39:67:@7311.16]
  wire [2:0] _GEN_21; // @[Conditional.scala 39:67:@7287.14]
  wire [2:0] _GEN_22; // @[Conditional.scala 39:67:@7248.12]
  wire [2:0] _GEN_23; // @[Conditional.scala 39:67:@7241.10]
  wire [2:0] _GEN_24; // @[Conditional.scala 39:67:@7234.8]
  wire [2:0] _GEN_25; // @[Conditional.scala 39:67:@7221.6]
  wire [2:0] _GEN_26; // @[Conditional.scala 40:58:@7203.4]
  wire  _T_640; // @[TensorLoad.scala 147:30:@7317.4]
  wire  _T_641; // @[TensorLoad.scala 147:40:@7318.4]
  wire  _T_643; // @[Decoupled.scala 37:37:@7324.4]
  wire  _T_648; // @[TensorLoad.scala 156:36:@7334.6]
  wire  _GEN_27; // @[TensorLoad.scala 156:57:@7335.6]
  wire  _GEN_28; // @[TensorLoad.scala 154:25:@7329.4]
  wire  _T_653; // @[TensorLoad.scala 161:44:@7340.4]
  wire  _T_660; // @[TensorLoad.scala 164:61:@7346.4]
  wire  _T_661; // @[TensorLoad.scala 164:48:@7347.4]
  wire  _T_662; // @[TensorLoad.scala 165:14:@7348.4]
  wire  _T_663; // @[TensorLoad.scala 165:25:@7349.4]
  wire  _T_664; // @[TensorLoad.scala 165:45:@7350.4]
  wire  _T_665; // @[TensorLoad.scala 164:70:@7351.4]
  wire  _T_671; // @[TensorLoad.scala 169:14:@7357.4]
  wire  _T_672; // @[TensorLoad.scala 169:25:@7358.4]
  wire  _T_673; // @[TensorLoad.scala 168:35:@7359.4]
  wire  _T_675; // @[TensorLoad.scala 170:32:@7361.4]
  wire  _T_676; // @[TensorLoad.scala 170:30:@7362.4]
  wire  _T_677; // @[TensorLoad.scala 170:46:@7363.4]
  wire  _T_680; // @[TensorLoad.scala 170:67:@7365.4]
  wire  _T_681; // @[TensorLoad.scala 169:46:@7366.4]
  wire  _T_685; // @[TensorLoad.scala 171:45:@7370.4]
  wire  _T_686; // @[TensorLoad.scala 170:89:@7371.4]
  wire  _T_691; // @[TensorLoad.scala 173:44:@7376.4]
  wire  _T_692; // @[TensorLoad.scala 174:28:@7377.4]
  wire  _T_693; // @[TensorLoad.scala 174:46:@7378.4]
  wire  _T_696; // @[TensorLoad.scala 174:67:@7380.4]
  wire  _T_697; // @[TensorLoad.scala 174:25:@7381.4]
  wire  _T_699; // @[TensorLoad.scala 182:32:@7388.4]
  wire  _T_702; // @[TensorLoad.scala 190:11:@7395.4]
  wire  _T_703; // @[TensorLoad.scala 189:36:@7396.4]
  wire  _T_705; // @[TensorLoad.scala 190:22:@7398.4]
  wire  _T_706; // @[TensorLoad.scala 192:11:@7399.4]
  wire  isZeroPad; // @[TensorLoad.scala 191:22:@7400.4]
  wire  _T_709; // @[TensorLoad.scala 194:24:@7403.4]
  wire  _T_711; // @[TensorLoad.scala 194:53:@7404.4]
  wire  _T_712; // @[TensorLoad.scala 194:46:@7405.4]
  wire  _T_715; // @[TensorLoad.scala 196:36:@7411.6]
  wire [3:0] _T_717; // @[TensorLoad.scala 197:16:@7413.8]
  wire [2:0] _T_718; // @[TensorLoad.scala 197:16:@7414.8]
  wire [2:0] _GEN_29; // @[TensorLoad.scala 196:50:@7412.6]
  wire  _T_732; // @[TensorLoad.scala 202:51:@7430.6]
  reg [10:0] waddr_cur; // @[TensorLoad.scala 206:22:@7436.4]
  reg [31:0] _RAND_11;
  reg [10:0] waddr_nxt; // @[TensorLoad.scala 207:22:@7437.4]
  reg [31:0] _RAND_12;
  wire [11:0] _T_748; // @[TensorLoad.scala 215:28:@7451.8]
  wire [10:0] _T_749; // @[TensorLoad.scala 215:28:@7452.8]
  wire  _T_751; // @[TensorLoad.scala 216:33:@7457.8]
  wire [15:0] _GEN_126; // @[TensorLoad.scala 217:28:@7459.10]
  wire [16:0] _T_752; // @[TensorLoad.scala 217:28:@7459.10]
  wire [15:0] _T_753; // @[TensorLoad.scala 217:28:@7460.10]
  wire [15:0] _GEN_33; // @[TensorLoad.scala 216:59:@7458.8]
  wire [15:0] _GEN_34; // @[TensorLoad.scala 216:59:@7458.8]
  wire [15:0] _GEN_35; // @[TensorLoad.scala 214:3:@7450.6]
  wire [15:0] _GEN_36; // @[TensorLoad.scala 214:3:@7450.6]
  wire [15:0] _GEN_37; // @[TensorLoad.scala 208:25:@7439.4]
  wire [15:0] _GEN_38; // @[TensorLoad.scala 208:25:@7439.4]
  wire  wmask_0_0; // @[TensorLoad.scala 235:26:@7478.4]
  wire [63:0] wdata_0_0; // @[TensorLoad.scala 236:25:@7480.4]
  wire  wmask_0_1; // @[TensorLoad.scala 235:26:@7482.4]
  wire  wmask_0_2; // @[TensorLoad.scala 235:26:@7486.4]
  wire  wmask_0_3; // @[TensorLoad.scala 235:26:@7490.4]
  wire  wmask_0_4; // @[TensorLoad.scala 235:26:@7494.4]
  wire  wmask_0_5; // @[TensorLoad.scala 235:26:@7498.4]
  wire  wmask_0_6; // @[TensorLoad.scala 235:26:@7502.4]
  wire [255:0] _T_855; // @[TensorLoad.scala 238:43:@7516.4]
  wire [511:0] _T_863; // @[TensorLoad.scala 238:43:@7524.4]
  wire [63:0] _T_915; // @[TensorLoad.scala 238:58:@7528.4]
  wire [63:0] _T_916; // @[TensorLoad.scala 238:58:@7530.4]
  wire [63:0] _T_917; // @[TensorLoad.scala 238:58:@7532.4]
  wire [63:0] _T_918; // @[TensorLoad.scala 238:58:@7534.4]
  wire [63:0] _T_919; // @[TensorLoad.scala 238:58:@7536.4]
  wire [63:0] _T_920; // @[TensorLoad.scala 238:58:@7538.4]
  wire [63:0] _T_921; // @[TensorLoad.scala 238:58:@7540.4]
  wire [63:0] _T_922; // @[TensorLoad.scala 238:58:@7542.4]
  reg  rvalid; // @[TensorLoad.scala 252:23:@7583.4]
  reg [31:0] _RAND_13;
  wire  _GEN_75; // @[TensorLoad.scala 256:26:@7588.4]
  wire [511:0] _T_1043; // @[TensorLoad.scala 259:38:@7600.4]
  wire  _T_1191; // @[TensorLoad.scala 263:96:@7656.4]
  wire  done_no_pad; // @[TensorLoad.scala 263:83:@7657.4]
  wire  done_x_pad; // @[TensorLoad.scala 264:72:@7662.4]
  wire  _T_1198; // @[TensorLoad.scala 265:37:@7664.4]
  wire  done_y_pad; // @[TensorLoad.scala 265:52:@7665.4]
  wire  _T_1199; // @[TensorLoad.scala 266:26:@7666.4]
  reg [10:0] tensorFile_0_0_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [10:0] tensorFile_0_1_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [10:0] tensorFile_0_2_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_16;
  reg [10:0] tensorFile_0_3_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [10:0] tensorFile_0_4_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_18;
  reg [10:0] tensorFile_0_5_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [10:0] tensorFile_0_6_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_20;
  reg [10:0] tensorFile_0_7_rdata_0_addr_pipe_0;
  reg [31:0] _RAND_21;
  TensorDataCtrl_2 dataCtrl ( // @[TensorLoad.scala 52:24:@7183.4]
    .clock(dataCtrl_clock),
    .io_start(dataCtrl_io_start),
    .io_done(dataCtrl_io_done),
    .io_inst(dataCtrl_io_inst),
    .io_baddr(dataCtrl_io_baddr),
    .io_xinit(dataCtrl_io_xinit),
    .io_xupdate(dataCtrl_io_xupdate),
    .io_yupdate(dataCtrl_io_yupdate),
    .io_stride(dataCtrl_io_stride),
    .io_split(dataCtrl_io_split),
    .io_addr(dataCtrl_io_addr),
    .io_len(dataCtrl_io_len)
  );
  TensorPadCtrl_8 yPadCtrl0 ( // @[TensorLoad.scala 55:25:@7187.4]
    .clock(yPadCtrl0_clock),
    .reset(yPadCtrl0_reset),
    .io_start(yPadCtrl0_io_start),
    .io_done(yPadCtrl0_io_done),
    .io_inst(yPadCtrl0_io_inst)
  );
  TensorPadCtrl_9 yPadCtrl1 ( // @[TensorLoad.scala 56:25:@7190.4]
    .clock(yPadCtrl1_clock),
    .reset(yPadCtrl1_reset),
    .io_start(yPadCtrl1_io_start),
    .io_done(yPadCtrl1_io_done),
    .io_inst(yPadCtrl1_io_inst)
  );
  TensorPadCtrl_10 xPadCtrl0 ( // @[TensorLoad.scala 57:25:@7193.4]
    .clock(xPadCtrl0_clock),
    .reset(xPadCtrl0_reset),
    .io_start(xPadCtrl0_io_start),
    .io_done(xPadCtrl0_io_done),
    .io_inst(xPadCtrl0_io_inst)
  );
  TensorPadCtrl_11 xPadCtrl1 ( // @[TensorLoad.scala 58:25:@7196.4]
    .clock(xPadCtrl1_clock),
    .reset(xPadCtrl1_reset),
    .io_start(xPadCtrl1_io_start),
    .io_done(xPadCtrl1_io_done),
    .io_inst(xPadCtrl1_io_inst)
  );
  assign tensorFile_0_0_rdata_0_addr = tensorFile_0_0_rdata_0_addr_pipe_0;
  assign tensorFile_0_0_rdata_0_data = tensorFile_0_0[tensorFile_0_0_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7466.4]
  assign tensorFile_0_0__T_992_data = _T_640 ? _T_915 : wdata_0_0;
  assign tensorFile_0_0__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_0__T_992_mask = _T_640 ? 1'h1 : wmask_0_0;
  assign tensorFile_0_0__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_1_rdata_0_addr = tensorFile_0_1_rdata_0_addr_pipe_0;
  assign tensorFile_0_1_rdata_0_data = tensorFile_0_1[tensorFile_0_1_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7466.4]
  assign tensorFile_0_1__T_992_data = _T_640 ? _T_916 : wdata_0_0;
  assign tensorFile_0_1__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_1__T_992_mask = _T_640 ? 1'h1 : wmask_0_1;
  assign tensorFile_0_1__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_2_rdata_0_addr = tensorFile_0_2_rdata_0_addr_pipe_0;
  assign tensorFile_0_2_rdata_0_data = tensorFile_0_2[tensorFile_0_2_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7466.4]
  assign tensorFile_0_2__T_992_data = _T_640 ? _T_917 : wdata_0_0;
  assign tensorFile_0_2__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_2__T_992_mask = _T_640 ? 1'h1 : wmask_0_2;
  assign tensorFile_0_2__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_3_rdata_0_addr = tensorFile_0_3_rdata_0_addr_pipe_0;
  assign tensorFile_0_3_rdata_0_data = tensorFile_0_3[tensorFile_0_3_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7466.4]
  assign tensorFile_0_3__T_992_data = _T_640 ? _T_918 : wdata_0_0;
  assign tensorFile_0_3__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_3__T_992_mask = _T_640 ? 1'h1 : wmask_0_3;
  assign tensorFile_0_3__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_4_rdata_0_addr = tensorFile_0_4_rdata_0_addr_pipe_0;
  assign tensorFile_0_4_rdata_0_data = tensorFile_0_4[tensorFile_0_4_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7466.4]
  assign tensorFile_0_4__T_992_data = _T_640 ? _T_919 : wdata_0_0;
  assign tensorFile_0_4__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_4__T_992_mask = _T_640 ? 1'h1 : wmask_0_4;
  assign tensorFile_0_4__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_5_rdata_0_addr = tensorFile_0_5_rdata_0_addr_pipe_0;
  assign tensorFile_0_5_rdata_0_data = tensorFile_0_5[tensorFile_0_5_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7466.4]
  assign tensorFile_0_5__T_992_data = _T_640 ? _T_920 : wdata_0_0;
  assign tensorFile_0_5__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_5__T_992_mask = _T_640 ? 1'h1 : wmask_0_5;
  assign tensorFile_0_5__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_6_rdata_0_addr = tensorFile_0_6_rdata_0_addr_pipe_0;
  assign tensorFile_0_6_rdata_0_data = tensorFile_0_6[tensorFile_0_6_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7466.4]
  assign tensorFile_0_6__T_992_data = _T_640 ? _T_921 : wdata_0_0;
  assign tensorFile_0_6__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_6__T_992_mask = _T_640 ? 1'h1 : wmask_0_6;
  assign tensorFile_0_6__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign tensorFile_0_7_rdata_0_addr = tensorFile_0_7_rdata_0_addr_pipe_0;
  assign tensorFile_0_7_rdata_0_data = tensorFile_0_7[tensorFile_0_7_rdata_0_addr]; // @[TensorLoad.scala 222:16:@7466.4]
  assign tensorFile_0_7__T_992_data = _T_640 ? _T_922 : wdata_0_0;
  assign tensorFile_0_7__T_992_addr = _T_640 ? io_tensor_wr_bits_idx : waddr_cur;
  assign tensorFile_0_7__T_992_mask = _T_640 ? 1'h1 : _T_711;
  assign tensorFile_0_7__T_992_en = _T_640 ? io_tensor_wr_valid : _T_715;
  assign dec_sram_offset = io_inst[24:9]; // @[TensorLoad.scala 51:29:@7163.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorLoad.scala 51:29:@7171.4]
  assign dec_ypad_0 = io_inst[115:112]; // @[TensorLoad.scala 51:29:@7175.4]
  assign dec_ypad_1 = io_inst[119:116]; // @[TensorLoad.scala 51:29:@7177.4]
  assign dec_xpad_0 = io_inst[123:120]; // @[TensorLoad.scala 51:29:@7179.4]
  assign dec_xpad_1 = io_inst[127:124]; // @[TensorLoad.scala 51:29:@7181.4]
  assign _T_614 = 3'h0 == state; // @[Conditional.scala 37:30:@7202.4]
  assign _T_616 = dec_ypad_0 != 4'h0; // @[TensorLoad.scala 71:25:@7205.8]
  assign _T_618 = dec_xpad_0 != 4'h0; // @[TensorLoad.scala 73:31:@7210.10]
  assign _GEN_0 = _T_618 ? 3'h2 : 3'h3; // @[TensorLoad.scala 73:40:@7211.10]
  assign _GEN_1 = _T_616 ? 3'h1 : _GEN_0; // @[TensorLoad.scala 71:34:@7206.8]
  assign _GEN_2 = io_start ? _GEN_1 : state; // @[TensorLoad.scala 70:22:@7204.6]
  assign _T_619 = 3'h1 == state; // @[Conditional.scala 37:30:@7220.6]
  assign _GEN_4 = yPadCtrl0_io_done ? _GEN_0 : state; // @[TensorLoad.scala 81:31:@7222.8]
  assign _T_622 = 3'h2 == state; // @[Conditional.scala 37:30:@7233.8]
  assign _GEN_5 = xPadCtrl0_io_done ? 3'h3 : state; // @[TensorLoad.scala 90:31:@7235.10]
  assign _T_623 = 3'h3 == state; // @[Conditional.scala 37:30:@7240.10]
  assign _GEN_6 = io_vme_rd_cmd_ready ? 3'h4 : state; // @[TensorLoad.scala 95:33:@7242.12]
  assign _T_624 = 3'h4 == state; // @[Conditional.scala 37:30:@7247.12]
  assign _T_626 = dec_xpad_1 != 4'h0; // @[TensorLoad.scala 102:27:@7251.18]
  assign _T_628 = dec_ypad_1 != 4'h0; // @[TensorLoad.scala 104:33:@7256.20]
  assign _GEN_7 = _T_628 ? 3'h6 : 3'h0; // @[TensorLoad.scala 104:42:@7257.20]
  assign _GEN_8 = _T_626 ? 3'h5 : _GEN_7; // @[TensorLoad.scala 102:36:@7252.18]
  assign _GEN_10 = _T_626 ? 3'h5 : _GEN_0; // @[TensorLoad.scala 110:36:@7267.20]
  assign _GEN_11 = dataCtrl_io_split ? 3'h3 : state; // @[TensorLoad.scala 117:39:@7280.20]
  assign _GEN_12 = dataCtrl_io_stride ? _GEN_10 : _GEN_11; // @[TensorLoad.scala 109:40:@7265.18]
  assign _GEN_13 = dataCtrl_io_done ? _GEN_8 : _GEN_12; // @[TensorLoad.scala 101:32:@7250.16]
  assign _GEN_14 = io_vme_rd_data_valid ? _GEN_13 : state; // @[TensorLoad.scala 100:34:@7249.14]
  assign _T_633 = 3'h5 == state; // @[Conditional.scala 37:30:@7286.14]
  assign _GEN_17 = dataCtrlDone ? _GEN_7 : _GEN_0; // @[TensorLoad.scala 124:28:@7289.18]
  assign _GEN_18 = xPadCtrl1_io_done ? _GEN_17 : state; // @[TensorLoad.scala 123:31:@7288.16]
  assign _T_638 = 3'h6 == state; // @[Conditional.scala 37:30:@7310.16]
  assign _T_639 = yPadCtrl1_io_done & dataCtrlDone; // @[TensorLoad.scala 140:30:@7312.18]
  assign _GEN_19 = _T_639 ? 3'h0 : state; // @[TensorLoad.scala 140:47:@7313.18]
  assign _GEN_20 = _T_638 ? _GEN_19 : state; // @[Conditional.scala 39:67:@7311.16]
  assign _GEN_21 = _T_633 ? _GEN_18 : _GEN_20; // @[Conditional.scala 39:67:@7287.14]
  assign _GEN_22 = _T_624 ? _GEN_14 : _GEN_21; // @[Conditional.scala 39:67:@7248.12]
  assign _GEN_23 = _T_623 ? _GEN_6 : _GEN_22; // @[Conditional.scala 39:67:@7241.10]
  assign _GEN_24 = _T_622 ? _GEN_5 : _GEN_23; // @[Conditional.scala 39:67:@7234.8]
  assign _GEN_25 = _T_619 ? _GEN_4 : _GEN_24; // @[Conditional.scala 39:67:@7221.6]
  assign _GEN_26 = _T_614 ? _GEN_2 : _GEN_25; // @[Conditional.scala 40:58:@7203.4]
  assign _T_640 = state == 3'h0; // @[TensorLoad.scala 147:30:@7317.4]
  assign _T_641 = _T_640 & io_start; // @[TensorLoad.scala 147:40:@7318.4]
  assign _T_643 = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[Decoupled.scala 37:37:@7324.4]
  assign _T_648 = _T_643 & dataCtrl_io_done; // @[TensorLoad.scala 156:36:@7334.6]
  assign _GEN_27 = _T_648 ? 1'h1 : dataCtrlDone; // @[TensorLoad.scala 156:57:@7335.6]
  assign _GEN_28 = _T_640 ? 1'h0 : _GEN_27; // @[TensorLoad.scala 154:25:@7329.4]
  assign _T_653 = _T_616 & _T_640; // @[TensorLoad.scala 161:44:@7340.4]
  assign _T_660 = dec_xpad_1 == 4'h0; // @[TensorLoad.scala 164:61:@7346.4]
  assign _T_661 = _T_648 & _T_660; // @[TensorLoad.scala 164:48:@7347.4]
  assign _T_662 = state == 3'h5; // @[TensorLoad.scala 165:14:@7348.4]
  assign _T_663 = _T_662 & xPadCtrl1_io_done; // @[TensorLoad.scala 165:25:@7349.4]
  assign _T_664 = _T_663 & dataCtrlDone; // @[TensorLoad.scala 165:45:@7350.4]
  assign _T_665 = _T_661 | _T_664; // @[TensorLoad.scala 164:70:@7351.4]
  assign _T_671 = state == 3'h1; // @[TensorLoad.scala 169:14:@7357.4]
  assign _T_672 = _T_671 & yPadCtrl0_io_done; // @[TensorLoad.scala 169:25:@7358.4]
  assign _T_673 = _T_641 | _T_672; // @[TensorLoad.scala 168:35:@7359.4]
  assign _T_675 = ~ dataCtrlDone; // @[TensorLoad.scala 170:32:@7361.4]
  assign _T_676 = _T_643 & _T_675; // @[TensorLoad.scala 170:30:@7362.4]
  assign _T_677 = _T_676 & dataCtrl_io_stride; // @[TensorLoad.scala 170:46:@7363.4]
  assign _T_680 = _T_677 & _T_660; // @[TensorLoad.scala 170:67:@7365.4]
  assign _T_681 = _T_673 | _T_680; // @[TensorLoad.scala 169:46:@7366.4]
  assign _T_685 = _T_663 & _T_675; // @[TensorLoad.scala 171:45:@7370.4]
  assign _T_686 = _T_681 | _T_685; // @[TensorLoad.scala 170:89:@7371.4]
  assign _T_691 = _T_626 & _T_643; // @[TensorLoad.scala 173:44:@7376.4]
  assign _T_692 = ~ dataCtrl_io_done; // @[TensorLoad.scala 174:28:@7377.4]
  assign _T_693 = _T_692 & dataCtrl_io_stride; // @[TensorLoad.scala 174:46:@7378.4]
  assign _T_696 = _T_693 & _T_626; // @[TensorLoad.scala 174:67:@7380.4]
  assign _T_697 = dataCtrl_io_done | _T_696; // @[TensorLoad.scala 174:25:@7381.4]
  assign _T_699 = state == 3'h3; // @[TensorLoad.scala 182:32:@7388.4]
  assign _T_702 = state == 3'h2; // @[TensorLoad.scala 190:11:@7395.4]
  assign _T_703 = _T_671 | _T_702; // @[TensorLoad.scala 189:36:@7396.4]
  assign _T_705 = _T_703 | _T_662; // @[TensorLoad.scala 190:22:@7398.4]
  assign _T_706 = state == 3'h6; // @[TensorLoad.scala 192:11:@7399.4]
  assign isZeroPad = _T_705 | _T_706; // @[TensorLoad.scala 191:22:@7400.4]
  assign _T_709 = _T_640 | _T_699; // @[TensorLoad.scala 194:24:@7403.4]
  assign _T_711 = tag == 3'h7; // @[TensorLoad.scala 194:53:@7404.4]
  assign _T_712 = _T_709 | _T_711; // @[TensorLoad.scala 194:46:@7405.4]
  assign _T_715 = _T_643 | isZeroPad; // @[TensorLoad.scala 196:36:@7411.6]
  assign _T_717 = tag + 3'h1; // @[TensorLoad.scala 197:16:@7413.8]
  assign _T_718 = tag + 3'h1; // @[TensorLoad.scala 197:16:@7414.8]
  assign _GEN_29 = _T_715 ? _T_718 : tag; // @[TensorLoad.scala 196:50:@7412.6]
  assign _T_732 = _T_715 & _T_711; // @[TensorLoad.scala 202:51:@7430.6]
  assign _T_748 = waddr_cur + 11'h1; // @[TensorLoad.scala 215:28:@7451.8]
  assign _T_749 = waddr_cur + 11'h1; // @[TensorLoad.scala 215:28:@7452.8]
  assign _T_751 = dataCtrl_io_stride & _T_643; // @[TensorLoad.scala 216:33:@7457.8]
  assign _GEN_126 = {{5'd0}, waddr_nxt}; // @[TensorLoad.scala 217:28:@7459.10]
  assign _T_752 = _GEN_126 + dec_xsize; // @[TensorLoad.scala 217:28:@7459.10]
  assign _T_753 = _GEN_126 + dec_xsize; // @[TensorLoad.scala 217:28:@7460.10]
  assign _GEN_33 = _T_751 ? _T_753 : {{5'd0}, waddr_cur}; // @[TensorLoad.scala 216:59:@7458.8]
  assign _GEN_34 = _T_751 ? _T_753 : {{5'd0}, waddr_nxt}; // @[TensorLoad.scala 216:59:@7458.8]
  assign _GEN_35 = _T_732 ? {{5'd0}, _T_749} : _GEN_33; // @[TensorLoad.scala 214:3:@7450.6]
  assign _GEN_36 = _T_732 ? {{5'd0}, waddr_nxt} : _GEN_34; // @[TensorLoad.scala 214:3:@7450.6]
  assign _GEN_37 = _T_640 ? dec_sram_offset : _GEN_35; // @[TensorLoad.scala 208:25:@7439.4]
  assign _GEN_38 = _T_640 ? dec_sram_offset : _GEN_36; // @[TensorLoad.scala 208:25:@7439.4]
  assign wmask_0_0 = tag == 3'h0; // @[TensorLoad.scala 235:26:@7478.4]
  assign wdata_0_0 = isZeroPad ? 64'h0 : io_vme_rd_data_bits; // @[TensorLoad.scala 236:25:@7480.4]
  assign wmask_0_1 = tag == 3'h1; // @[TensorLoad.scala 235:26:@7482.4]
  assign wmask_0_2 = tag == 3'h2; // @[TensorLoad.scala 235:26:@7486.4]
  assign wmask_0_3 = tag == 3'h3; // @[TensorLoad.scala 235:26:@7490.4]
  assign wmask_0_4 = tag == 3'h4; // @[TensorLoad.scala 235:26:@7494.4]
  assign wmask_0_5 = tag == 3'h5; // @[TensorLoad.scala 235:26:@7498.4]
  assign wmask_0_6 = tag == 3'h6; // @[TensorLoad.scala 235:26:@7502.4]
  assign _T_855 = {io_tensor_wr_bits_data_0_7,io_tensor_wr_bits_data_0_6,io_tensor_wr_bits_data_0_5,io_tensor_wr_bits_data_0_4,io_tensor_wr_bits_data_0_3,io_tensor_wr_bits_data_0_2,io_tensor_wr_bits_data_0_1,io_tensor_wr_bits_data_0_0}; // @[TensorLoad.scala 238:43:@7516.4]
  assign _T_863 = {io_tensor_wr_bits_data_0_15,io_tensor_wr_bits_data_0_14,io_tensor_wr_bits_data_0_13,io_tensor_wr_bits_data_0_12,io_tensor_wr_bits_data_0_11,io_tensor_wr_bits_data_0_10,io_tensor_wr_bits_data_0_9,io_tensor_wr_bits_data_0_8,_T_855}; // @[TensorLoad.scala 238:43:@7524.4]
  assign _T_915 = _T_863[63:0]; // @[TensorLoad.scala 238:58:@7528.4]
  assign _T_916 = _T_863[127:64]; // @[TensorLoad.scala 238:58:@7530.4]
  assign _T_917 = _T_863[191:128]; // @[TensorLoad.scala 238:58:@7532.4]
  assign _T_918 = _T_863[255:192]; // @[TensorLoad.scala 238:58:@7534.4]
  assign _T_919 = _T_863[319:256]; // @[TensorLoad.scala 238:58:@7536.4]
  assign _T_920 = _T_863[383:320]; // @[TensorLoad.scala 238:58:@7538.4]
  assign _T_921 = _T_863[447:384]; // @[TensorLoad.scala 238:58:@7540.4]
  assign _T_922 = _T_863[511:448]; // @[TensorLoad.scala 238:58:@7542.4]
  assign _GEN_75 = io_tensor_rd_idx_valid; // @[TensorLoad.scala 256:26:@7588.4]
  assign _T_1043 = {tensorFile_0_7_rdata_0_data,tensorFile_0_6_rdata_0_data,tensorFile_0_5_rdata_0_data,tensorFile_0_4_rdata_0_data,tensorFile_0_3_rdata_0_data,tensorFile_0_2_rdata_0_data,tensorFile_0_1_rdata_0_data,tensorFile_0_0_rdata_0_data}; // @[TensorLoad.scala 259:38:@7600.4]
  assign _T_1191 = dec_ypad_1 == 4'h0; // @[TensorLoad.scala 263:96:@7656.4]
  assign done_no_pad = _T_661 & _T_1191; // @[TensorLoad.scala 263:83:@7657.4]
  assign done_x_pad = _T_664 & _T_1191; // @[TensorLoad.scala 264:72:@7662.4]
  assign _T_1198 = _T_706 & dataCtrlDone; // @[TensorLoad.scala 265:37:@7664.4]
  assign done_y_pad = _T_1198 & yPadCtrl1_io_done; // @[TensorLoad.scala 265:52:@7665.4]
  assign _T_1199 = done_no_pad | done_x_pad; // @[TensorLoad.scala 266:26:@7666.4]
  assign io_done = _T_1199 | done_y_pad; // @[TensorLoad.scala 266:11:@7668.4]
  assign io_vme_rd_cmd_valid = state == 3'h3; // @[TensorLoad.scala 182:23:@7389.4]
  assign io_vme_rd_cmd_bits_addr = dataCtrl_io_addr; // @[TensorLoad.scala 183:27:@7390.4]
  assign io_vme_rd_cmd_bits_len = dataCtrl_io_len; // @[TensorLoad.scala 184:26:@7391.4]
  assign io_vme_rd_data_ready = state == 3'h4; // @[TensorLoad.scala 186:24:@7393.4]
  assign io_tensor_rd_data_valid = rvalid; // @[TensorLoad.scala 253:27:@7585.4]
  assign io_tensor_rd_data_bits_0_0 = _T_1043[31:0]; // @[TensorLoad.scala 259:33:@7636.4]
  assign io_tensor_rd_data_bits_0_1 = _T_1043[63:32]; // @[TensorLoad.scala 259:33:@7637.4]
  assign io_tensor_rd_data_bits_0_2 = _T_1043[95:64]; // @[TensorLoad.scala 259:33:@7638.4]
  assign io_tensor_rd_data_bits_0_3 = _T_1043[127:96]; // @[TensorLoad.scala 259:33:@7639.4]
  assign io_tensor_rd_data_bits_0_4 = _T_1043[159:128]; // @[TensorLoad.scala 259:33:@7640.4]
  assign io_tensor_rd_data_bits_0_5 = _T_1043[191:160]; // @[TensorLoad.scala 259:33:@7641.4]
  assign io_tensor_rd_data_bits_0_6 = _T_1043[223:192]; // @[TensorLoad.scala 259:33:@7642.4]
  assign io_tensor_rd_data_bits_0_7 = _T_1043[255:224]; // @[TensorLoad.scala 259:33:@7643.4]
  assign io_tensor_rd_data_bits_0_8 = _T_1043[287:256]; // @[TensorLoad.scala 259:33:@7644.4]
  assign io_tensor_rd_data_bits_0_9 = _T_1043[319:288]; // @[TensorLoad.scala 259:33:@7645.4]
  assign io_tensor_rd_data_bits_0_10 = _T_1043[351:320]; // @[TensorLoad.scala 259:33:@7646.4]
  assign io_tensor_rd_data_bits_0_11 = _T_1043[383:352]; // @[TensorLoad.scala 259:33:@7647.4]
  assign io_tensor_rd_data_bits_0_12 = _T_1043[415:384]; // @[TensorLoad.scala 259:33:@7648.4]
  assign io_tensor_rd_data_bits_0_13 = _T_1043[447:416]; // @[TensorLoad.scala 259:33:@7649.4]
  assign io_tensor_rd_data_bits_0_14 = _T_1043[479:448]; // @[TensorLoad.scala 259:33:@7650.4]
  assign io_tensor_rd_data_bits_0_15 = _T_1043[511:480]; // @[TensorLoad.scala 259:33:@7651.4]
  assign dataCtrl_clock = clock; // @[:@7184.4]
  assign dataCtrl_io_start = _T_640 & io_start; // @[TensorLoad.scala 147:21:@7319.4]
  assign dataCtrl_io_inst = io_inst; // @[TensorLoad.scala 148:20:@7320.4]
  assign dataCtrl_io_baddr = io_baddr; // @[TensorLoad.scala 149:21:@7321.4]
  assign dataCtrl_io_xinit = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[TensorLoad.scala 150:21:@7323.4]
  assign dataCtrl_io_xupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 151:23:@7325.4]
  assign dataCtrl_io_yupdate = io_vme_rd_data_ready & io_vme_rd_data_valid; // @[TensorLoad.scala 152:23:@7327.4]
  assign yPadCtrl0_clock = clock; // @[:@7188.4]
  assign yPadCtrl0_reset = reset; // @[:@7189.4]
  assign yPadCtrl0_io_start = _T_653 & io_start; // @[TensorLoad.scala 161:22:@7342.4]
  assign yPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 176:21:@7384.4]
  assign yPadCtrl1_clock = clock; // @[:@7191.4]
  assign yPadCtrl1_reset = reset; // @[:@7192.4]
  assign yPadCtrl1_io_start = _T_628 & _T_665; // @[TensorLoad.scala 163:22:@7353.4]
  assign yPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 177:21:@7385.4]
  assign xPadCtrl0_clock = clock; // @[:@7194.4]
  assign xPadCtrl0_reset = reset; // @[:@7195.4]
  assign xPadCtrl0_io_start = _T_618 & _T_686; // @[TensorLoad.scala 167:22:@7373.4]
  assign xPadCtrl0_io_inst = io_inst; // @[TensorLoad.scala 178:21:@7386.4]
  assign xPadCtrl1_clock = clock; // @[:@7197.4]
  assign xPadCtrl1_reset = reset; // @[:@7198.4]
  assign xPadCtrl1_io_start = _T_691 & _T_697; // @[TensorLoad.scala 173:22:@7383.4]
  assign xPadCtrl1_io_inst = io_inst; // @[TensorLoad.scala 179:21:@7387.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_0[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_1[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_2[initvar] = _RAND_2[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_3[initvar] = _RAND_3[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_4[initvar] = _RAND_4[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_5[initvar] = _RAND_5[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_6[initvar] = _RAND_6[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_7[initvar] = _RAND_7[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  dataCtrlDone = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  tag = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  waddr_cur = _RAND_11[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  waddr_nxt = _RAND_12[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  rvalid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  tensorFile_0_0_rdata_0_addr_pipe_0 = _RAND_14[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  tensorFile_0_1_rdata_0_addr_pipe_0 = _RAND_15[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  tensorFile_0_2_rdata_0_addr_pipe_0 = _RAND_16[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  tensorFile_0_3_rdata_0_addr_pipe_0 = _RAND_17[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  tensorFile_0_4_rdata_0_addr_pipe_0 = _RAND_18[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  tensorFile_0_5_rdata_0_addr_pipe_0 = _RAND_19[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  tensorFile_0_6_rdata_0_addr_pipe_0 = _RAND_20[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  tensorFile_0_7_rdata_0_addr_pipe_0 = _RAND_21[10:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tensorFile_0_0__T_992_en & tensorFile_0_0__T_992_mask) begin
      tensorFile_0_0[tensorFile_0_0__T_992_addr] <= tensorFile_0_0__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
    end
    if(tensorFile_0_1__T_992_en & tensorFile_0_1__T_992_mask) begin
      tensorFile_0_1[tensorFile_0_1__T_992_addr] <= tensorFile_0_1__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
    end
    if(tensorFile_0_2__T_992_en & tensorFile_0_2__T_992_mask) begin
      tensorFile_0_2[tensorFile_0_2__T_992_addr] <= tensorFile_0_2__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
    end
    if(tensorFile_0_3__T_992_en & tensorFile_0_3__T_992_mask) begin
      tensorFile_0_3[tensorFile_0_3__T_992_addr] <= tensorFile_0_3__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
    end
    if(tensorFile_0_4__T_992_en & tensorFile_0_4__T_992_mask) begin
      tensorFile_0_4[tensorFile_0_4__T_992_addr] <= tensorFile_0_4__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
    end
    if(tensorFile_0_5__T_992_en & tensorFile_0_5__T_992_mask) begin
      tensorFile_0_5[tensorFile_0_5__T_992_addr] <= tensorFile_0_5__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
    end
    if(tensorFile_0_6__T_992_en & tensorFile_0_6__T_992_mask) begin
      tensorFile_0_6[tensorFile_0_6__T_992_addr] <= tensorFile_0_6__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
    end
    if(tensorFile_0_7__T_992_en & tensorFile_0_7__T_992_mask) begin
      tensorFile_0_7[tensorFile_0_7__T_992_addr] <= tensorFile_0_7__T_992_data; // @[TensorLoad.scala 222:16:@7466.4]
    end
    if (reset) begin
      dataCtrlDone <= 1'h0;
    end else begin
      if (_T_640) begin
        dataCtrlDone <= 1'h0;
      end else begin
        if (_T_648) begin
          dataCtrlDone <= 1'h1;
        end
      end
    end
    if (_T_712) begin
      tag <= 3'h0;
    end else begin
      if (_T_715) begin
        tag <= _T_718;
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_614) begin
        if (io_start) begin
          if (_T_616) begin
            state <= 3'h1;
          end else begin
            if (_T_618) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end
      end else begin
        if (_T_619) begin
          if (yPadCtrl0_io_done) begin
            if (_T_618) begin
              state <= 3'h2;
            end else begin
              state <= 3'h3;
            end
          end
        end else begin
          if (_T_622) begin
            if (xPadCtrl0_io_done) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_623) begin
              if (io_vme_rd_cmd_ready) begin
                state <= 3'h4;
              end
            end else begin
              if (_T_624) begin
                if (io_vme_rd_data_valid) begin
                  if (dataCtrl_io_done) begin
                    if (_T_626) begin
                      state <= 3'h5;
                    end else begin
                      if (_T_628) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end
                  end else begin
                    if (dataCtrl_io_stride) begin
                      if (_T_626) begin
                        state <= 3'h5;
                      end else begin
                        if (_T_618) begin
                          state <= 3'h2;
                        end else begin
                          state <= 3'h3;
                        end
                      end
                    end else begin
                      if (dataCtrl_io_split) begin
                        state <= 3'h3;
                      end
                    end
                  end
                end
              end else begin
                if (_T_633) begin
                  if (xPadCtrl1_io_done) begin
                    if (dataCtrlDone) begin
                      if (_T_628) begin
                        state <= 3'h6;
                      end else begin
                        state <= 3'h0;
                      end
                    end else begin
                      if (_T_618) begin
                        state <= 3'h2;
                      end else begin
                        state <= 3'h3;
                      end
                    end
                  end
                end else begin
                  if (_T_638) begin
                    if (_T_639) begin
                      state <= 3'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    waddr_cur <= _GEN_37[10:0];
    waddr_nxt <= _GEN_38[10:0];
    rvalid <= io_tensor_rd_idx_valid;
    if (_GEN_75) begin
      tensorFile_0_0_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_1_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_2_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_3_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_4_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_5_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_6_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
    if (_GEN_75) begin
      tensorFile_0_7_rdata_0_addr_pipe_0 <= io_tensor_rd_idx_bits;
    end
  end
endmodule
module MAC( // @[:@7670.2]
  input         clock, // @[:@7671.4]
  input  [7:0]  io_a, // @[:@7673.4]
  input  [7:0]  io_b, // @[:@7673.4]
  input         io_c, // @[:@7673.4]
  output [16:0] io_y // @[:@7673.4]
);
  reg [7:0] rA; // @[TensorGemm.scala 39:19:@7677.4]
  reg [31:0] _RAND_0;
  reg [7:0] rB; // @[TensorGemm.scala 40:19:@7679.4]
  reg [31:0] _RAND_1;
  reg  rC; // @[TensorGemm.scala 41:19:@7681.4]
  reg [31:0] _RAND_2;
  wire [15:0] mult; // @[TensorGemm.scala 43:14:@7683.4]
  wire [15:0] _GEN_0; // @[TensorGemm.scala 44:13:@7685.4]
  assign mult = $signed(rA) * $signed(rB); // @[TensorGemm.scala 43:14:@7683.4]
  assign _GEN_0 = {16{rC}}; // @[TensorGemm.scala 44:13:@7685.4]
  assign io_y = $signed(_GEN_0) + $signed(mult); // @[TensorGemm.scala 46:8:@7687.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rA = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rB = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rC = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    rA <= io_a;
    rB <= io_b;
    rC <= io_c;
  end
endmodule
module PipeAdder( // @[:@7974.2]
  input         clock, // @[:@7975.4]
  input  [16:0] io_a, // @[:@7977.4]
  input  [16:0] io_b, // @[:@7977.4]
  output [17:0] io_y // @[:@7977.4]
);
  reg [16:0] rA; // @[TensorGemm.scala 61:19:@7980.4]
  reg [31:0] _RAND_0;
  reg [16:0] rB; // @[TensorGemm.scala 62:19:@7982.4]
  reg [31:0] _RAND_1;
  assign io_y = $signed(rA) + $signed(rB); // @[TensorGemm.scala 64:8:@7986.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rA = _RAND_0[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rB = _RAND_1[16:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    rA <= io_a;
    rB <= io_b;
  end
endmodule
module Adder( // @[:@8086.2]
  input  [17:0] io_a, // @[:@8089.4]
  input  [17:0] io_b, // @[:@8089.4]
  output [18:0] io_y // @[:@8089.4]
);
  assign io_y = $signed(io_a) + $signed(io_b); // @[TensorGemm.scala 85:8:@8098.4]
endmodule
module Adder_4( // @[:@8142.2]
  input  [18:0] io_a, // @[:@8145.4]
  input  [18:0] io_b, // @[:@8145.4]
  output [19:0] io_y // @[:@8145.4]
);
  assign io_y = $signed(io_a) + $signed(io_b); // @[TensorGemm.scala 85:8:@8154.4]
endmodule
module Adder_6( // @[:@8170.2]
  input  [19:0] io_a, // @[:@8173.4]
  input  [19:0] io_b, // @[:@8173.4]
  output [20:0] io_y // @[:@8173.4]
);
  assign io_y = $signed(io_a) + $signed(io_b); // @[TensorGemm.scala 85:8:@8182.4]
endmodule
module DotProduct( // @[:@8184.2]
  input         clock, // @[:@8185.4]
  input  [7:0]  io_a_0, // @[:@8187.4]
  input  [7:0]  io_a_1, // @[:@8187.4]
  input  [7:0]  io_a_2, // @[:@8187.4]
  input  [7:0]  io_a_3, // @[:@8187.4]
  input  [7:0]  io_a_4, // @[:@8187.4]
  input  [7:0]  io_a_5, // @[:@8187.4]
  input  [7:0]  io_a_6, // @[:@8187.4]
  input  [7:0]  io_a_7, // @[:@8187.4]
  input  [7:0]  io_a_8, // @[:@8187.4]
  input  [7:0]  io_a_9, // @[:@8187.4]
  input  [7:0]  io_a_10, // @[:@8187.4]
  input  [7:0]  io_a_11, // @[:@8187.4]
  input  [7:0]  io_a_12, // @[:@8187.4]
  input  [7:0]  io_a_13, // @[:@8187.4]
  input  [7:0]  io_a_14, // @[:@8187.4]
  input  [7:0]  io_a_15, // @[:@8187.4]
  input  [7:0]  io_b_0, // @[:@8187.4]
  input  [7:0]  io_b_1, // @[:@8187.4]
  input  [7:0]  io_b_2, // @[:@8187.4]
  input  [7:0]  io_b_3, // @[:@8187.4]
  input  [7:0]  io_b_4, // @[:@8187.4]
  input  [7:0]  io_b_5, // @[:@8187.4]
  input  [7:0]  io_b_6, // @[:@8187.4]
  input  [7:0]  io_b_7, // @[:@8187.4]
  input  [7:0]  io_b_8, // @[:@8187.4]
  input  [7:0]  io_b_9, // @[:@8187.4]
  input  [7:0]  io_b_10, // @[:@8187.4]
  input  [7:0]  io_b_11, // @[:@8187.4]
  input  [7:0]  io_b_12, // @[:@8187.4]
  input  [7:0]  io_b_13, // @[:@8187.4]
  input  [7:0]  io_b_14, // @[:@8187.4]
  input  [7:0]  io_b_15, // @[:@8187.4]
  output [20:0] io_y // @[:@8187.4]
);
  wire  m_0_clock; // @[TensorGemm.scala 103:32:@8189.4]
  wire [7:0] m_0_io_a; // @[TensorGemm.scala 103:32:@8189.4]
  wire [7:0] m_0_io_b; // @[TensorGemm.scala 103:32:@8189.4]
  wire  m_0_io_c; // @[TensorGemm.scala 103:32:@8189.4]
  wire [16:0] m_0_io_y; // @[TensorGemm.scala 103:32:@8189.4]
  wire  m_1_clock; // @[TensorGemm.scala 103:32:@8192.4]
  wire [7:0] m_1_io_a; // @[TensorGemm.scala 103:32:@8192.4]
  wire [7:0] m_1_io_b; // @[TensorGemm.scala 103:32:@8192.4]
  wire  m_1_io_c; // @[TensorGemm.scala 103:32:@8192.4]
  wire [16:0] m_1_io_y; // @[TensorGemm.scala 103:32:@8192.4]
  wire  m_2_clock; // @[TensorGemm.scala 103:32:@8195.4]
  wire [7:0] m_2_io_a; // @[TensorGemm.scala 103:32:@8195.4]
  wire [7:0] m_2_io_b; // @[TensorGemm.scala 103:32:@8195.4]
  wire  m_2_io_c; // @[TensorGemm.scala 103:32:@8195.4]
  wire [16:0] m_2_io_y; // @[TensorGemm.scala 103:32:@8195.4]
  wire  m_3_clock; // @[TensorGemm.scala 103:32:@8198.4]
  wire [7:0] m_3_io_a; // @[TensorGemm.scala 103:32:@8198.4]
  wire [7:0] m_3_io_b; // @[TensorGemm.scala 103:32:@8198.4]
  wire  m_3_io_c; // @[TensorGemm.scala 103:32:@8198.4]
  wire [16:0] m_3_io_y; // @[TensorGemm.scala 103:32:@8198.4]
  wire  m_4_clock; // @[TensorGemm.scala 103:32:@8201.4]
  wire [7:0] m_4_io_a; // @[TensorGemm.scala 103:32:@8201.4]
  wire [7:0] m_4_io_b; // @[TensorGemm.scala 103:32:@8201.4]
  wire  m_4_io_c; // @[TensorGemm.scala 103:32:@8201.4]
  wire [16:0] m_4_io_y; // @[TensorGemm.scala 103:32:@8201.4]
  wire  m_5_clock; // @[TensorGemm.scala 103:32:@8204.4]
  wire [7:0] m_5_io_a; // @[TensorGemm.scala 103:32:@8204.4]
  wire [7:0] m_5_io_b; // @[TensorGemm.scala 103:32:@8204.4]
  wire  m_5_io_c; // @[TensorGemm.scala 103:32:@8204.4]
  wire [16:0] m_5_io_y; // @[TensorGemm.scala 103:32:@8204.4]
  wire  m_6_clock; // @[TensorGemm.scala 103:32:@8207.4]
  wire [7:0] m_6_io_a; // @[TensorGemm.scala 103:32:@8207.4]
  wire [7:0] m_6_io_b; // @[TensorGemm.scala 103:32:@8207.4]
  wire  m_6_io_c; // @[TensorGemm.scala 103:32:@8207.4]
  wire [16:0] m_6_io_y; // @[TensorGemm.scala 103:32:@8207.4]
  wire  m_7_clock; // @[TensorGemm.scala 103:32:@8210.4]
  wire [7:0] m_7_io_a; // @[TensorGemm.scala 103:32:@8210.4]
  wire [7:0] m_7_io_b; // @[TensorGemm.scala 103:32:@8210.4]
  wire  m_7_io_c; // @[TensorGemm.scala 103:32:@8210.4]
  wire [16:0] m_7_io_y; // @[TensorGemm.scala 103:32:@8210.4]
  wire  m_8_clock; // @[TensorGemm.scala 103:32:@8213.4]
  wire [7:0] m_8_io_a; // @[TensorGemm.scala 103:32:@8213.4]
  wire [7:0] m_8_io_b; // @[TensorGemm.scala 103:32:@8213.4]
  wire  m_8_io_c; // @[TensorGemm.scala 103:32:@8213.4]
  wire [16:0] m_8_io_y; // @[TensorGemm.scala 103:32:@8213.4]
  wire  m_9_clock; // @[TensorGemm.scala 103:32:@8216.4]
  wire [7:0] m_9_io_a; // @[TensorGemm.scala 103:32:@8216.4]
  wire [7:0] m_9_io_b; // @[TensorGemm.scala 103:32:@8216.4]
  wire  m_9_io_c; // @[TensorGemm.scala 103:32:@8216.4]
  wire [16:0] m_9_io_y; // @[TensorGemm.scala 103:32:@8216.4]
  wire  m_10_clock; // @[TensorGemm.scala 103:32:@8219.4]
  wire [7:0] m_10_io_a; // @[TensorGemm.scala 103:32:@8219.4]
  wire [7:0] m_10_io_b; // @[TensorGemm.scala 103:32:@8219.4]
  wire  m_10_io_c; // @[TensorGemm.scala 103:32:@8219.4]
  wire [16:0] m_10_io_y; // @[TensorGemm.scala 103:32:@8219.4]
  wire  m_11_clock; // @[TensorGemm.scala 103:32:@8222.4]
  wire [7:0] m_11_io_a; // @[TensorGemm.scala 103:32:@8222.4]
  wire [7:0] m_11_io_b; // @[TensorGemm.scala 103:32:@8222.4]
  wire  m_11_io_c; // @[TensorGemm.scala 103:32:@8222.4]
  wire [16:0] m_11_io_y; // @[TensorGemm.scala 103:32:@8222.4]
  wire  m_12_clock; // @[TensorGemm.scala 103:32:@8225.4]
  wire [7:0] m_12_io_a; // @[TensorGemm.scala 103:32:@8225.4]
  wire [7:0] m_12_io_b; // @[TensorGemm.scala 103:32:@8225.4]
  wire  m_12_io_c; // @[TensorGemm.scala 103:32:@8225.4]
  wire [16:0] m_12_io_y; // @[TensorGemm.scala 103:32:@8225.4]
  wire  m_13_clock; // @[TensorGemm.scala 103:32:@8228.4]
  wire [7:0] m_13_io_a; // @[TensorGemm.scala 103:32:@8228.4]
  wire [7:0] m_13_io_b; // @[TensorGemm.scala 103:32:@8228.4]
  wire  m_13_io_c; // @[TensorGemm.scala 103:32:@8228.4]
  wire [16:0] m_13_io_y; // @[TensorGemm.scala 103:32:@8228.4]
  wire  m_14_clock; // @[TensorGemm.scala 103:32:@8231.4]
  wire [7:0] m_14_io_a; // @[TensorGemm.scala 103:32:@8231.4]
  wire [7:0] m_14_io_b; // @[TensorGemm.scala 103:32:@8231.4]
  wire  m_14_io_c; // @[TensorGemm.scala 103:32:@8231.4]
  wire [16:0] m_14_io_y; // @[TensorGemm.scala 103:32:@8231.4]
  wire  m_15_clock; // @[TensorGemm.scala 103:32:@8234.4]
  wire [7:0] m_15_io_a; // @[TensorGemm.scala 103:32:@8234.4]
  wire [7:0] m_15_io_b; // @[TensorGemm.scala 103:32:@8234.4]
  wire  m_15_io_c; // @[TensorGemm.scala 103:32:@8234.4]
  wire [16:0] m_15_io_y; // @[TensorGemm.scala 103:32:@8234.4]
  wire  a_0_0_clock; // @[TensorGemm.scala 108:17:@8237.4]
  wire [16:0] a_0_0_io_a; // @[TensorGemm.scala 108:17:@8237.4]
  wire [16:0] a_0_0_io_b; // @[TensorGemm.scala 108:17:@8237.4]
  wire [17:0] a_0_0_io_y; // @[TensorGemm.scala 108:17:@8237.4]
  wire  a_0_1_clock; // @[TensorGemm.scala 108:17:@8240.4]
  wire [16:0] a_0_1_io_a; // @[TensorGemm.scala 108:17:@8240.4]
  wire [16:0] a_0_1_io_b; // @[TensorGemm.scala 108:17:@8240.4]
  wire [17:0] a_0_1_io_y; // @[TensorGemm.scala 108:17:@8240.4]
  wire  a_0_2_clock; // @[TensorGemm.scala 108:17:@8243.4]
  wire [16:0] a_0_2_io_a; // @[TensorGemm.scala 108:17:@8243.4]
  wire [16:0] a_0_2_io_b; // @[TensorGemm.scala 108:17:@8243.4]
  wire [17:0] a_0_2_io_y; // @[TensorGemm.scala 108:17:@8243.4]
  wire  a_0_3_clock; // @[TensorGemm.scala 108:17:@8246.4]
  wire [16:0] a_0_3_io_a; // @[TensorGemm.scala 108:17:@8246.4]
  wire [16:0] a_0_3_io_b; // @[TensorGemm.scala 108:17:@8246.4]
  wire [17:0] a_0_3_io_y; // @[TensorGemm.scala 108:17:@8246.4]
  wire  a_0_4_clock; // @[TensorGemm.scala 108:17:@8249.4]
  wire [16:0] a_0_4_io_a; // @[TensorGemm.scala 108:17:@8249.4]
  wire [16:0] a_0_4_io_b; // @[TensorGemm.scala 108:17:@8249.4]
  wire [17:0] a_0_4_io_y; // @[TensorGemm.scala 108:17:@8249.4]
  wire  a_0_5_clock; // @[TensorGemm.scala 108:17:@8252.4]
  wire [16:0] a_0_5_io_a; // @[TensorGemm.scala 108:17:@8252.4]
  wire [16:0] a_0_5_io_b; // @[TensorGemm.scala 108:17:@8252.4]
  wire [17:0] a_0_5_io_y; // @[TensorGemm.scala 108:17:@8252.4]
  wire  a_0_6_clock; // @[TensorGemm.scala 108:17:@8255.4]
  wire [16:0] a_0_6_io_a; // @[TensorGemm.scala 108:17:@8255.4]
  wire [16:0] a_0_6_io_b; // @[TensorGemm.scala 108:17:@8255.4]
  wire [17:0] a_0_6_io_y; // @[TensorGemm.scala 108:17:@8255.4]
  wire  a_0_7_clock; // @[TensorGemm.scala 108:17:@8258.4]
  wire [16:0] a_0_7_io_a; // @[TensorGemm.scala 108:17:@8258.4]
  wire [16:0] a_0_7_io_b; // @[TensorGemm.scala 108:17:@8258.4]
  wire [17:0] a_0_7_io_y; // @[TensorGemm.scala 108:17:@8258.4]
  wire [17:0] a_1_0_io_a; // @[TensorGemm.scala 110:17:@8261.4]
  wire [17:0] a_1_0_io_b; // @[TensorGemm.scala 110:17:@8261.4]
  wire [18:0] a_1_0_io_y; // @[TensorGemm.scala 110:17:@8261.4]
  wire [17:0] a_1_1_io_a; // @[TensorGemm.scala 110:17:@8264.4]
  wire [17:0] a_1_1_io_b; // @[TensorGemm.scala 110:17:@8264.4]
  wire [18:0] a_1_1_io_y; // @[TensorGemm.scala 110:17:@8264.4]
  wire [17:0] a_1_2_io_a; // @[TensorGemm.scala 110:17:@8267.4]
  wire [17:0] a_1_2_io_b; // @[TensorGemm.scala 110:17:@8267.4]
  wire [18:0] a_1_2_io_y; // @[TensorGemm.scala 110:17:@8267.4]
  wire [17:0] a_1_3_io_a; // @[TensorGemm.scala 110:17:@8270.4]
  wire [17:0] a_1_3_io_b; // @[TensorGemm.scala 110:17:@8270.4]
  wire [18:0] a_1_3_io_y; // @[TensorGemm.scala 110:17:@8270.4]
  wire [18:0] a_2_0_io_a; // @[TensorGemm.scala 110:17:@8273.4]
  wire [18:0] a_2_0_io_b; // @[TensorGemm.scala 110:17:@8273.4]
  wire [19:0] a_2_0_io_y; // @[TensorGemm.scala 110:17:@8273.4]
  wire [18:0] a_2_1_io_a; // @[TensorGemm.scala 110:17:@8276.4]
  wire [18:0] a_2_1_io_b; // @[TensorGemm.scala 110:17:@8276.4]
  wire [19:0] a_2_1_io_y; // @[TensorGemm.scala 110:17:@8276.4]
  wire [19:0] a_3_0_io_a; // @[TensorGemm.scala 110:17:@8279.4]
  wire [19:0] a_3_0_io_b; // @[TensorGemm.scala 110:17:@8279.4]
  wire [20:0] a_3_0_io_y; // @[TensorGemm.scala 110:17:@8279.4]
  MAC m_0 ( // @[TensorGemm.scala 103:32:@8189.4]
    .clock(m_0_clock),
    .io_a(m_0_io_a),
    .io_b(m_0_io_b),
    .io_c(m_0_io_c),
    .io_y(m_0_io_y)
  );
  MAC m_1 ( // @[TensorGemm.scala 103:32:@8192.4]
    .clock(m_1_clock),
    .io_a(m_1_io_a),
    .io_b(m_1_io_b),
    .io_c(m_1_io_c),
    .io_y(m_1_io_y)
  );
  MAC m_2 ( // @[TensorGemm.scala 103:32:@8195.4]
    .clock(m_2_clock),
    .io_a(m_2_io_a),
    .io_b(m_2_io_b),
    .io_c(m_2_io_c),
    .io_y(m_2_io_y)
  );
  MAC m_3 ( // @[TensorGemm.scala 103:32:@8198.4]
    .clock(m_3_clock),
    .io_a(m_3_io_a),
    .io_b(m_3_io_b),
    .io_c(m_3_io_c),
    .io_y(m_3_io_y)
  );
  MAC m_4 ( // @[TensorGemm.scala 103:32:@8201.4]
    .clock(m_4_clock),
    .io_a(m_4_io_a),
    .io_b(m_4_io_b),
    .io_c(m_4_io_c),
    .io_y(m_4_io_y)
  );
  MAC m_5 ( // @[TensorGemm.scala 103:32:@8204.4]
    .clock(m_5_clock),
    .io_a(m_5_io_a),
    .io_b(m_5_io_b),
    .io_c(m_5_io_c),
    .io_y(m_5_io_y)
  );
  MAC m_6 ( // @[TensorGemm.scala 103:32:@8207.4]
    .clock(m_6_clock),
    .io_a(m_6_io_a),
    .io_b(m_6_io_b),
    .io_c(m_6_io_c),
    .io_y(m_6_io_y)
  );
  MAC m_7 ( // @[TensorGemm.scala 103:32:@8210.4]
    .clock(m_7_clock),
    .io_a(m_7_io_a),
    .io_b(m_7_io_b),
    .io_c(m_7_io_c),
    .io_y(m_7_io_y)
  );
  MAC m_8 ( // @[TensorGemm.scala 103:32:@8213.4]
    .clock(m_8_clock),
    .io_a(m_8_io_a),
    .io_b(m_8_io_b),
    .io_c(m_8_io_c),
    .io_y(m_8_io_y)
  );
  MAC m_9 ( // @[TensorGemm.scala 103:32:@8216.4]
    .clock(m_9_clock),
    .io_a(m_9_io_a),
    .io_b(m_9_io_b),
    .io_c(m_9_io_c),
    .io_y(m_9_io_y)
  );
  MAC m_10 ( // @[TensorGemm.scala 103:32:@8219.4]
    .clock(m_10_clock),
    .io_a(m_10_io_a),
    .io_b(m_10_io_b),
    .io_c(m_10_io_c),
    .io_y(m_10_io_y)
  );
  MAC m_11 ( // @[TensorGemm.scala 103:32:@8222.4]
    .clock(m_11_clock),
    .io_a(m_11_io_a),
    .io_b(m_11_io_b),
    .io_c(m_11_io_c),
    .io_y(m_11_io_y)
  );
  MAC m_12 ( // @[TensorGemm.scala 103:32:@8225.4]
    .clock(m_12_clock),
    .io_a(m_12_io_a),
    .io_b(m_12_io_b),
    .io_c(m_12_io_c),
    .io_y(m_12_io_y)
  );
  MAC m_13 ( // @[TensorGemm.scala 103:32:@8228.4]
    .clock(m_13_clock),
    .io_a(m_13_io_a),
    .io_b(m_13_io_b),
    .io_c(m_13_io_c),
    .io_y(m_13_io_y)
  );
  MAC m_14 ( // @[TensorGemm.scala 103:32:@8231.4]
    .clock(m_14_clock),
    .io_a(m_14_io_a),
    .io_b(m_14_io_b),
    .io_c(m_14_io_c),
    .io_y(m_14_io_y)
  );
  MAC m_15 ( // @[TensorGemm.scala 103:32:@8234.4]
    .clock(m_15_clock),
    .io_a(m_15_io_a),
    .io_b(m_15_io_b),
    .io_c(m_15_io_c),
    .io_y(m_15_io_y)
  );
  PipeAdder a_0_0 ( // @[TensorGemm.scala 108:17:@8237.4]
    .clock(a_0_0_clock),
    .io_a(a_0_0_io_a),
    .io_b(a_0_0_io_b),
    .io_y(a_0_0_io_y)
  );
  PipeAdder a_0_1 ( // @[TensorGemm.scala 108:17:@8240.4]
    .clock(a_0_1_clock),
    .io_a(a_0_1_io_a),
    .io_b(a_0_1_io_b),
    .io_y(a_0_1_io_y)
  );
  PipeAdder a_0_2 ( // @[TensorGemm.scala 108:17:@8243.4]
    .clock(a_0_2_clock),
    .io_a(a_0_2_io_a),
    .io_b(a_0_2_io_b),
    .io_y(a_0_2_io_y)
  );
  PipeAdder a_0_3 ( // @[TensorGemm.scala 108:17:@8246.4]
    .clock(a_0_3_clock),
    .io_a(a_0_3_io_a),
    .io_b(a_0_3_io_b),
    .io_y(a_0_3_io_y)
  );
  PipeAdder a_0_4 ( // @[TensorGemm.scala 108:17:@8249.4]
    .clock(a_0_4_clock),
    .io_a(a_0_4_io_a),
    .io_b(a_0_4_io_b),
    .io_y(a_0_4_io_y)
  );
  PipeAdder a_0_5 ( // @[TensorGemm.scala 108:17:@8252.4]
    .clock(a_0_5_clock),
    .io_a(a_0_5_io_a),
    .io_b(a_0_5_io_b),
    .io_y(a_0_5_io_y)
  );
  PipeAdder a_0_6 ( // @[TensorGemm.scala 108:17:@8255.4]
    .clock(a_0_6_clock),
    .io_a(a_0_6_io_a),
    .io_b(a_0_6_io_b),
    .io_y(a_0_6_io_y)
  );
  PipeAdder a_0_7 ( // @[TensorGemm.scala 108:17:@8258.4]
    .clock(a_0_7_clock),
    .io_a(a_0_7_io_a),
    .io_b(a_0_7_io_b),
    .io_y(a_0_7_io_y)
  );
  Adder a_1_0 ( // @[TensorGemm.scala 110:17:@8261.4]
    .io_a(a_1_0_io_a),
    .io_b(a_1_0_io_b),
    .io_y(a_1_0_io_y)
  );
  Adder a_1_1 ( // @[TensorGemm.scala 110:17:@8264.4]
    .io_a(a_1_1_io_a),
    .io_b(a_1_1_io_b),
    .io_y(a_1_1_io_y)
  );
  Adder a_1_2 ( // @[TensorGemm.scala 110:17:@8267.4]
    .io_a(a_1_2_io_a),
    .io_b(a_1_2_io_b),
    .io_y(a_1_2_io_y)
  );
  Adder a_1_3 ( // @[TensorGemm.scala 110:17:@8270.4]
    .io_a(a_1_3_io_a),
    .io_b(a_1_3_io_b),
    .io_y(a_1_3_io_y)
  );
  Adder_4 a_2_0 ( // @[TensorGemm.scala 110:17:@8273.4]
    .io_a(a_2_0_io_a),
    .io_b(a_2_0_io_b),
    .io_y(a_2_0_io_y)
  );
  Adder_4 a_2_1 ( // @[TensorGemm.scala 110:17:@8276.4]
    .io_a(a_2_1_io_a),
    .io_b(a_2_1_io_b),
    .io_y(a_2_1_io_y)
  );
  Adder_6 a_3_0 ( // @[TensorGemm.scala 110:17:@8279.4]
    .io_a(a_3_0_io_a),
    .io_b(a_3_0_io_b),
    .io_y(a_3_0_io_y)
  );
  assign io_y = a_3_0_io_y; // @[TensorGemm.scala 134:8:@8360.4]
  assign m_0_clock = clock; // @[:@8190.4]
  assign m_0_io_a = io_a_0; // @[TensorGemm.scala 114:15:@8282.4]
  assign m_0_io_b = io_b_0; // @[TensorGemm.scala 115:15:@8283.4]
  assign m_0_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8284.4]
  assign m_1_clock = clock; // @[:@8193.4]
  assign m_1_io_a = io_a_1; // @[TensorGemm.scala 114:15:@8285.4]
  assign m_1_io_b = io_b_1; // @[TensorGemm.scala 115:15:@8286.4]
  assign m_1_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8287.4]
  assign m_2_clock = clock; // @[:@8196.4]
  assign m_2_io_a = io_a_2; // @[TensorGemm.scala 114:15:@8288.4]
  assign m_2_io_b = io_b_2; // @[TensorGemm.scala 115:15:@8289.4]
  assign m_2_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8290.4]
  assign m_3_clock = clock; // @[:@8199.4]
  assign m_3_io_a = io_a_3; // @[TensorGemm.scala 114:15:@8291.4]
  assign m_3_io_b = io_b_3; // @[TensorGemm.scala 115:15:@8292.4]
  assign m_3_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8293.4]
  assign m_4_clock = clock; // @[:@8202.4]
  assign m_4_io_a = io_a_4; // @[TensorGemm.scala 114:15:@8294.4]
  assign m_4_io_b = io_b_4; // @[TensorGemm.scala 115:15:@8295.4]
  assign m_4_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8296.4]
  assign m_5_clock = clock; // @[:@8205.4]
  assign m_5_io_a = io_a_5; // @[TensorGemm.scala 114:15:@8297.4]
  assign m_5_io_b = io_b_5; // @[TensorGemm.scala 115:15:@8298.4]
  assign m_5_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8299.4]
  assign m_6_clock = clock; // @[:@8208.4]
  assign m_6_io_a = io_a_6; // @[TensorGemm.scala 114:15:@8300.4]
  assign m_6_io_b = io_b_6; // @[TensorGemm.scala 115:15:@8301.4]
  assign m_6_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8302.4]
  assign m_7_clock = clock; // @[:@8211.4]
  assign m_7_io_a = io_a_7; // @[TensorGemm.scala 114:15:@8303.4]
  assign m_7_io_b = io_b_7; // @[TensorGemm.scala 115:15:@8304.4]
  assign m_7_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8305.4]
  assign m_8_clock = clock; // @[:@8214.4]
  assign m_8_io_a = io_a_8; // @[TensorGemm.scala 114:15:@8306.4]
  assign m_8_io_b = io_b_8; // @[TensorGemm.scala 115:15:@8307.4]
  assign m_8_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8308.4]
  assign m_9_clock = clock; // @[:@8217.4]
  assign m_9_io_a = io_a_9; // @[TensorGemm.scala 114:15:@8309.4]
  assign m_9_io_b = io_b_9; // @[TensorGemm.scala 115:15:@8310.4]
  assign m_9_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8311.4]
  assign m_10_clock = clock; // @[:@8220.4]
  assign m_10_io_a = io_a_10; // @[TensorGemm.scala 114:15:@8312.4]
  assign m_10_io_b = io_b_10; // @[TensorGemm.scala 115:15:@8313.4]
  assign m_10_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8314.4]
  assign m_11_clock = clock; // @[:@8223.4]
  assign m_11_io_a = io_a_11; // @[TensorGemm.scala 114:15:@8315.4]
  assign m_11_io_b = io_b_11; // @[TensorGemm.scala 115:15:@8316.4]
  assign m_11_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8317.4]
  assign m_12_clock = clock; // @[:@8226.4]
  assign m_12_io_a = io_a_12; // @[TensorGemm.scala 114:15:@8318.4]
  assign m_12_io_b = io_b_12; // @[TensorGemm.scala 115:15:@8319.4]
  assign m_12_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8320.4]
  assign m_13_clock = clock; // @[:@8229.4]
  assign m_13_io_a = io_a_13; // @[TensorGemm.scala 114:15:@8321.4]
  assign m_13_io_b = io_b_13; // @[TensorGemm.scala 115:15:@8322.4]
  assign m_13_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8323.4]
  assign m_14_clock = clock; // @[:@8232.4]
  assign m_14_io_a = io_a_14; // @[TensorGemm.scala 114:15:@8324.4]
  assign m_14_io_b = io_b_14; // @[TensorGemm.scala 115:15:@8325.4]
  assign m_14_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8326.4]
  assign m_15_clock = clock; // @[:@8235.4]
  assign m_15_io_a = io_a_15; // @[TensorGemm.scala 114:15:@8327.4]
  assign m_15_io_b = io_b_15; // @[TensorGemm.scala 115:15:@8328.4]
  assign m_15_io_c = 1'sh0; // @[TensorGemm.scala 116:15:@8329.4]
  assign a_0_0_clock = clock; // @[:@8238.4]
  assign a_0_0_io_a = m_0_io_y; // @[TensorGemm.scala 124:22:@8330.4]
  assign a_0_0_io_b = m_1_io_y; // @[TensorGemm.scala 125:22:@8331.4]
  assign a_0_1_clock = clock; // @[:@8241.4]
  assign a_0_1_io_a = m_2_io_y; // @[TensorGemm.scala 124:22:@8332.4]
  assign a_0_1_io_b = m_3_io_y; // @[TensorGemm.scala 125:22:@8333.4]
  assign a_0_2_clock = clock; // @[:@8244.4]
  assign a_0_2_io_a = m_4_io_y; // @[TensorGemm.scala 124:22:@8334.4]
  assign a_0_2_io_b = m_5_io_y; // @[TensorGemm.scala 125:22:@8335.4]
  assign a_0_3_clock = clock; // @[:@8247.4]
  assign a_0_3_io_a = m_6_io_y; // @[TensorGemm.scala 124:22:@8336.4]
  assign a_0_3_io_b = m_7_io_y; // @[TensorGemm.scala 125:22:@8337.4]
  assign a_0_4_clock = clock; // @[:@8250.4]
  assign a_0_4_io_a = m_8_io_y; // @[TensorGemm.scala 124:22:@8338.4]
  assign a_0_4_io_b = m_9_io_y; // @[TensorGemm.scala 125:22:@8339.4]
  assign a_0_5_clock = clock; // @[:@8253.4]
  assign a_0_5_io_a = m_10_io_y; // @[TensorGemm.scala 124:22:@8340.4]
  assign a_0_5_io_b = m_11_io_y; // @[TensorGemm.scala 125:22:@8341.4]
  assign a_0_6_clock = clock; // @[:@8256.4]
  assign a_0_6_io_a = m_12_io_y; // @[TensorGemm.scala 124:22:@8342.4]
  assign a_0_6_io_b = m_13_io_y; // @[TensorGemm.scala 125:22:@8343.4]
  assign a_0_7_clock = clock; // @[:@8259.4]
  assign a_0_7_io_a = m_14_io_y; // @[TensorGemm.scala 124:22:@8344.4]
  assign a_0_7_io_b = m_15_io_y; // @[TensorGemm.scala 125:22:@8345.4]
  assign a_1_0_io_a = a_0_0_io_y; // @[TensorGemm.scala 127:22:@8346.4]
  assign a_1_0_io_b = a_0_1_io_y; // @[TensorGemm.scala 128:22:@8347.4]
  assign a_1_1_io_a = a_0_2_io_y; // @[TensorGemm.scala 127:22:@8348.4]
  assign a_1_1_io_b = a_0_3_io_y; // @[TensorGemm.scala 128:22:@8349.4]
  assign a_1_2_io_a = a_0_4_io_y; // @[TensorGemm.scala 127:22:@8350.4]
  assign a_1_2_io_b = a_0_5_io_y; // @[TensorGemm.scala 128:22:@8351.4]
  assign a_1_3_io_a = a_0_6_io_y; // @[TensorGemm.scala 127:22:@8352.4]
  assign a_1_3_io_b = a_0_7_io_y; // @[TensorGemm.scala 128:22:@8353.4]
  assign a_2_0_io_a = a_1_0_io_y; // @[TensorGemm.scala 127:22:@8354.4]
  assign a_2_0_io_b = a_1_1_io_y; // @[TensorGemm.scala 128:22:@8355.4]
  assign a_2_1_io_a = a_1_2_io_y; // @[TensorGemm.scala 127:22:@8356.4]
  assign a_2_1_io_b = a_1_3_io_y; // @[TensorGemm.scala 128:22:@8357.4]
  assign a_3_0_io_a = a_2_0_io_y; // @[TensorGemm.scala 127:22:@8358.4]
  assign a_3_0_io_b = a_2_1_io_y; // @[TensorGemm.scala 128:22:@8359.4]
endmodule
module Pipe( // @[:@18742.2]
  input         clock, // @[:@18743.4]
  input         reset, // @[:@18744.4]
  input         io_enq_valid, // @[:@18745.4]
  input  [31:0] io_enq_bits, // @[:@18745.4]
  output        io_deq_valid, // @[:@18745.4]
  output [31:0] io_deq_bits // @[:@18745.4]
);
  reg  _T_19; // @[Valid.scala 48:22:@18747.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_21; // @[Reg.scala 11:16:@18749.4]
  reg [31:0] _RAND_1;
  reg  _T_24; // @[Valid.scala 48:22:@18753.4]
  reg [31:0] _RAND_2;
  reg [31:0] _T_26; // @[Reg.scala 11:16:@18755.4]
  reg [31:0] _RAND_3;
  assign io_deq_valid = _T_24; // @[Valid.scala 70:10:@18763.4]
  assign io_deq_bits = _T_26; // @[Valid.scala 70:10:@18762.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_21 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_24 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_26 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      _T_19 <= io_enq_valid;
    end
    if (io_enq_valid) begin
      _T_21 <= io_enq_bits;
    end
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_19;
    end
    if (_T_19) begin
      _T_26 <= _T_21;
    end
  end
endmodule
module MatrixVectorMultiplication( // @[:@19110.2]
  input         clock, // @[:@19111.4]
  input         reset, // @[:@19112.4]
  input         io_reset, // @[:@19113.4]
  input         io_inp_data_valid, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_0, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_1, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_2, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_3, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_4, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_5, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_6, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_7, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_8, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_9, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_10, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_11, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_12, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_13, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_14, // @[:@19113.4]
  input  [7:0]  io_inp_data_bits_0_15, // @[:@19113.4]
  input         io_wgt_data_valid, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_0_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_1_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_2_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_3_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_4_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_5_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_6_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_7_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_8_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_9_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_10_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_11_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_12_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_13_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_14_15, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_0, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_1, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_2, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_3, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_4, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_5, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_6, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_7, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_8, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_9, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_10, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_11, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_12, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_13, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_14, // @[:@19113.4]
  input  [7:0]  io_wgt_data_bits_15_15, // @[:@19113.4]
  input         io_acc_i_data_valid, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_0, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_1, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_2, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_3, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_4, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_5, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_6, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_7, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_8, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_9, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_10, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_11, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_12, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_13, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_14, // @[:@19113.4]
  input  [31:0] io_acc_i_data_bits_0_15, // @[:@19113.4]
  output        io_acc_o_data_valid, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_0, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_1, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_2, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_3, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_4, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_5, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_6, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_7, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_8, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_9, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_10, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_11, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_12, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_13, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_14, // @[:@19113.4]
  output [31:0] io_acc_o_data_bits_0_15, // @[:@19113.4]
  output        io_out_data_valid, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_0, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_1, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_2, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_3, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_4, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_5, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_6, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_7, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_8, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_9, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_10, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_11, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_12, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_13, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_14, // @[:@19113.4]
  output [7:0]  io_out_data_bits_0_15 // @[:@19113.4]
);
  wire  dot_0_clock; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_0; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_1; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_2; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_3; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_4; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_5; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_6; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_7; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_8; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_9; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_10; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_11; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_12; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_13; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_14; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_a_15; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_0; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_1; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_2; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_3; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_4; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_5; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_6; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_7; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_8; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_9; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_10; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_11; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_12; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_13; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_14; // @[TensorGemm.scala 153:11:@19115.4]
  wire [7:0] dot_0_io_b_15; // @[TensorGemm.scala 153:11:@19115.4]
  wire [20:0] dot_0_io_y; // @[TensorGemm.scala 153:11:@19115.4]
  wire  dot_1_clock; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_0; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_1; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_2; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_3; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_4; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_5; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_6; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_7; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_8; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_9; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_10; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_11; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_12; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_13; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_14; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_a_15; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_0; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_1; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_2; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_3; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_4; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_5; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_6; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_7; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_8; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_9; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_10; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_11; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_12; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_13; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_14; // @[TensorGemm.scala 153:11:@19118.4]
  wire [7:0] dot_1_io_b_15; // @[TensorGemm.scala 153:11:@19118.4]
  wire [20:0] dot_1_io_y; // @[TensorGemm.scala 153:11:@19118.4]
  wire  dot_2_clock; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_0; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_1; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_2; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_3; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_4; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_5; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_6; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_7; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_8; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_9; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_10; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_11; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_12; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_13; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_14; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_a_15; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_0; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_1; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_2; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_3; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_4; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_5; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_6; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_7; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_8; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_9; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_10; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_11; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_12; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_13; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_14; // @[TensorGemm.scala 153:11:@19121.4]
  wire [7:0] dot_2_io_b_15; // @[TensorGemm.scala 153:11:@19121.4]
  wire [20:0] dot_2_io_y; // @[TensorGemm.scala 153:11:@19121.4]
  wire  dot_3_clock; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_0; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_1; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_2; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_3; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_4; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_5; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_6; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_7; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_8; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_9; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_10; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_11; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_12; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_13; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_14; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_a_15; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_0; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_1; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_2; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_3; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_4; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_5; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_6; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_7; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_8; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_9; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_10; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_11; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_12; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_13; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_14; // @[TensorGemm.scala 153:11:@19124.4]
  wire [7:0] dot_3_io_b_15; // @[TensorGemm.scala 153:11:@19124.4]
  wire [20:0] dot_3_io_y; // @[TensorGemm.scala 153:11:@19124.4]
  wire  dot_4_clock; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_0; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_1; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_2; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_3; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_4; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_5; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_6; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_7; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_8; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_9; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_10; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_11; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_12; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_13; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_14; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_a_15; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_0; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_1; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_2; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_3; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_4; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_5; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_6; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_7; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_8; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_9; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_10; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_11; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_12; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_13; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_14; // @[TensorGemm.scala 153:11:@19127.4]
  wire [7:0] dot_4_io_b_15; // @[TensorGemm.scala 153:11:@19127.4]
  wire [20:0] dot_4_io_y; // @[TensorGemm.scala 153:11:@19127.4]
  wire  dot_5_clock; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_0; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_1; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_2; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_3; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_4; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_5; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_6; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_7; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_8; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_9; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_10; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_11; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_12; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_13; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_14; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_a_15; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_0; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_1; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_2; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_3; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_4; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_5; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_6; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_7; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_8; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_9; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_10; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_11; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_12; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_13; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_14; // @[TensorGemm.scala 153:11:@19130.4]
  wire [7:0] dot_5_io_b_15; // @[TensorGemm.scala 153:11:@19130.4]
  wire [20:0] dot_5_io_y; // @[TensorGemm.scala 153:11:@19130.4]
  wire  dot_6_clock; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_0; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_1; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_2; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_3; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_4; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_5; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_6; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_7; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_8; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_9; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_10; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_11; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_12; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_13; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_14; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_a_15; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_0; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_1; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_2; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_3; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_4; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_5; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_6; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_7; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_8; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_9; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_10; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_11; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_12; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_13; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_14; // @[TensorGemm.scala 153:11:@19133.4]
  wire [7:0] dot_6_io_b_15; // @[TensorGemm.scala 153:11:@19133.4]
  wire [20:0] dot_6_io_y; // @[TensorGemm.scala 153:11:@19133.4]
  wire  dot_7_clock; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_0; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_1; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_2; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_3; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_4; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_5; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_6; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_7; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_8; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_9; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_10; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_11; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_12; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_13; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_14; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_a_15; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_0; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_1; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_2; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_3; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_4; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_5; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_6; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_7; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_8; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_9; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_10; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_11; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_12; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_13; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_14; // @[TensorGemm.scala 153:11:@19136.4]
  wire [7:0] dot_7_io_b_15; // @[TensorGemm.scala 153:11:@19136.4]
  wire [20:0] dot_7_io_y; // @[TensorGemm.scala 153:11:@19136.4]
  wire  dot_8_clock; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_0; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_1; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_2; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_3; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_4; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_5; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_6; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_7; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_8; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_9; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_10; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_11; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_12; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_13; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_14; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_a_15; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_0; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_1; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_2; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_3; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_4; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_5; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_6; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_7; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_8; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_9; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_10; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_11; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_12; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_13; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_14; // @[TensorGemm.scala 153:11:@19139.4]
  wire [7:0] dot_8_io_b_15; // @[TensorGemm.scala 153:11:@19139.4]
  wire [20:0] dot_8_io_y; // @[TensorGemm.scala 153:11:@19139.4]
  wire  dot_9_clock; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_0; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_1; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_2; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_3; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_4; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_5; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_6; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_7; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_8; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_9; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_10; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_11; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_12; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_13; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_14; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_a_15; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_0; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_1; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_2; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_3; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_4; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_5; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_6; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_7; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_8; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_9; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_10; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_11; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_12; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_13; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_14; // @[TensorGemm.scala 153:11:@19142.4]
  wire [7:0] dot_9_io_b_15; // @[TensorGemm.scala 153:11:@19142.4]
  wire [20:0] dot_9_io_y; // @[TensorGemm.scala 153:11:@19142.4]
  wire  dot_10_clock; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_0; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_1; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_2; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_3; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_4; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_5; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_6; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_7; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_8; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_9; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_10; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_11; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_12; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_13; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_14; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_a_15; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_0; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_1; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_2; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_3; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_4; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_5; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_6; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_7; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_8; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_9; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_10; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_11; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_12; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_13; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_14; // @[TensorGemm.scala 153:11:@19145.4]
  wire [7:0] dot_10_io_b_15; // @[TensorGemm.scala 153:11:@19145.4]
  wire [20:0] dot_10_io_y; // @[TensorGemm.scala 153:11:@19145.4]
  wire  dot_11_clock; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_0; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_1; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_2; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_3; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_4; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_5; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_6; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_7; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_8; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_9; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_10; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_11; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_12; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_13; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_14; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_a_15; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_0; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_1; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_2; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_3; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_4; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_5; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_6; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_7; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_8; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_9; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_10; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_11; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_12; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_13; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_14; // @[TensorGemm.scala 153:11:@19148.4]
  wire [7:0] dot_11_io_b_15; // @[TensorGemm.scala 153:11:@19148.4]
  wire [20:0] dot_11_io_y; // @[TensorGemm.scala 153:11:@19148.4]
  wire  dot_12_clock; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_0; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_1; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_2; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_3; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_4; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_5; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_6; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_7; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_8; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_9; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_10; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_11; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_12; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_13; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_14; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_a_15; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_0; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_1; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_2; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_3; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_4; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_5; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_6; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_7; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_8; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_9; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_10; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_11; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_12; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_13; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_14; // @[TensorGemm.scala 153:11:@19151.4]
  wire [7:0] dot_12_io_b_15; // @[TensorGemm.scala 153:11:@19151.4]
  wire [20:0] dot_12_io_y; // @[TensorGemm.scala 153:11:@19151.4]
  wire  dot_13_clock; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_0; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_1; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_2; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_3; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_4; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_5; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_6; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_7; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_8; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_9; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_10; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_11; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_12; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_13; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_14; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_a_15; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_0; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_1; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_2; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_3; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_4; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_5; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_6; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_7; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_8; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_9; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_10; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_11; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_12; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_13; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_14; // @[TensorGemm.scala 153:11:@19154.4]
  wire [7:0] dot_13_io_b_15; // @[TensorGemm.scala 153:11:@19154.4]
  wire [20:0] dot_13_io_y; // @[TensorGemm.scala 153:11:@19154.4]
  wire  dot_14_clock; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_0; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_1; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_2; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_3; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_4; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_5; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_6; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_7; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_8; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_9; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_10; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_11; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_12; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_13; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_14; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_a_15; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_0; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_1; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_2; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_3; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_4; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_5; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_6; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_7; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_8; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_9; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_10; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_11; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_12; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_13; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_14; // @[TensorGemm.scala 153:11:@19157.4]
  wire [7:0] dot_14_io_b_15; // @[TensorGemm.scala 153:11:@19157.4]
  wire [20:0] dot_14_io_y; // @[TensorGemm.scala 153:11:@19157.4]
  wire  dot_15_clock; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_0; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_1; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_2; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_3; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_4; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_5; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_6; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_7; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_8; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_9; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_10; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_11; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_12; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_13; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_14; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_a_15; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_0; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_1; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_2; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_3; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_4; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_5; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_6; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_7; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_8; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_9; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_10; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_11; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_12; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_13; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_14; // @[TensorGemm.scala 153:11:@19160.4]
  wire [7:0] dot_15_io_b_15; // @[TensorGemm.scala 153:11:@19160.4]
  wire [20:0] dot_15_io_y; // @[TensorGemm.scala 153:11:@19160.4]
  wire  acc_0_clock; // @[TensorGemm.scala 156:34:@19163.4]
  wire  acc_0_reset; // @[TensorGemm.scala 156:34:@19163.4]
  wire  acc_0_io_enq_valid; // @[TensorGemm.scala 156:34:@19163.4]
  wire [31:0] acc_0_io_enq_bits; // @[TensorGemm.scala 156:34:@19163.4]
  wire  acc_0_io_deq_valid; // @[TensorGemm.scala 156:34:@19163.4]
  wire [31:0] acc_0_io_deq_bits; // @[TensorGemm.scala 156:34:@19163.4]
  wire  acc_1_clock; // @[TensorGemm.scala 156:34:@19166.4]
  wire  acc_1_reset; // @[TensorGemm.scala 156:34:@19166.4]
  wire  acc_1_io_enq_valid; // @[TensorGemm.scala 156:34:@19166.4]
  wire [31:0] acc_1_io_enq_bits; // @[TensorGemm.scala 156:34:@19166.4]
  wire  acc_1_io_deq_valid; // @[TensorGemm.scala 156:34:@19166.4]
  wire [31:0] acc_1_io_deq_bits; // @[TensorGemm.scala 156:34:@19166.4]
  wire  acc_2_clock; // @[TensorGemm.scala 156:34:@19169.4]
  wire  acc_2_reset; // @[TensorGemm.scala 156:34:@19169.4]
  wire  acc_2_io_enq_valid; // @[TensorGemm.scala 156:34:@19169.4]
  wire [31:0] acc_2_io_enq_bits; // @[TensorGemm.scala 156:34:@19169.4]
  wire  acc_2_io_deq_valid; // @[TensorGemm.scala 156:34:@19169.4]
  wire [31:0] acc_2_io_deq_bits; // @[TensorGemm.scala 156:34:@19169.4]
  wire  acc_3_clock; // @[TensorGemm.scala 156:34:@19172.4]
  wire  acc_3_reset; // @[TensorGemm.scala 156:34:@19172.4]
  wire  acc_3_io_enq_valid; // @[TensorGemm.scala 156:34:@19172.4]
  wire [31:0] acc_3_io_enq_bits; // @[TensorGemm.scala 156:34:@19172.4]
  wire  acc_3_io_deq_valid; // @[TensorGemm.scala 156:34:@19172.4]
  wire [31:0] acc_3_io_deq_bits; // @[TensorGemm.scala 156:34:@19172.4]
  wire  acc_4_clock; // @[TensorGemm.scala 156:34:@19175.4]
  wire  acc_4_reset; // @[TensorGemm.scala 156:34:@19175.4]
  wire  acc_4_io_enq_valid; // @[TensorGemm.scala 156:34:@19175.4]
  wire [31:0] acc_4_io_enq_bits; // @[TensorGemm.scala 156:34:@19175.4]
  wire  acc_4_io_deq_valid; // @[TensorGemm.scala 156:34:@19175.4]
  wire [31:0] acc_4_io_deq_bits; // @[TensorGemm.scala 156:34:@19175.4]
  wire  acc_5_clock; // @[TensorGemm.scala 156:34:@19178.4]
  wire  acc_5_reset; // @[TensorGemm.scala 156:34:@19178.4]
  wire  acc_5_io_enq_valid; // @[TensorGemm.scala 156:34:@19178.4]
  wire [31:0] acc_5_io_enq_bits; // @[TensorGemm.scala 156:34:@19178.4]
  wire  acc_5_io_deq_valid; // @[TensorGemm.scala 156:34:@19178.4]
  wire [31:0] acc_5_io_deq_bits; // @[TensorGemm.scala 156:34:@19178.4]
  wire  acc_6_clock; // @[TensorGemm.scala 156:34:@19181.4]
  wire  acc_6_reset; // @[TensorGemm.scala 156:34:@19181.4]
  wire  acc_6_io_enq_valid; // @[TensorGemm.scala 156:34:@19181.4]
  wire [31:0] acc_6_io_enq_bits; // @[TensorGemm.scala 156:34:@19181.4]
  wire  acc_6_io_deq_valid; // @[TensorGemm.scala 156:34:@19181.4]
  wire [31:0] acc_6_io_deq_bits; // @[TensorGemm.scala 156:34:@19181.4]
  wire  acc_7_clock; // @[TensorGemm.scala 156:34:@19184.4]
  wire  acc_7_reset; // @[TensorGemm.scala 156:34:@19184.4]
  wire  acc_7_io_enq_valid; // @[TensorGemm.scala 156:34:@19184.4]
  wire [31:0] acc_7_io_enq_bits; // @[TensorGemm.scala 156:34:@19184.4]
  wire  acc_7_io_deq_valid; // @[TensorGemm.scala 156:34:@19184.4]
  wire [31:0] acc_7_io_deq_bits; // @[TensorGemm.scala 156:34:@19184.4]
  wire  acc_8_clock; // @[TensorGemm.scala 156:34:@19187.4]
  wire  acc_8_reset; // @[TensorGemm.scala 156:34:@19187.4]
  wire  acc_8_io_enq_valid; // @[TensorGemm.scala 156:34:@19187.4]
  wire [31:0] acc_8_io_enq_bits; // @[TensorGemm.scala 156:34:@19187.4]
  wire  acc_8_io_deq_valid; // @[TensorGemm.scala 156:34:@19187.4]
  wire [31:0] acc_8_io_deq_bits; // @[TensorGemm.scala 156:34:@19187.4]
  wire  acc_9_clock; // @[TensorGemm.scala 156:34:@19190.4]
  wire  acc_9_reset; // @[TensorGemm.scala 156:34:@19190.4]
  wire  acc_9_io_enq_valid; // @[TensorGemm.scala 156:34:@19190.4]
  wire [31:0] acc_9_io_enq_bits; // @[TensorGemm.scala 156:34:@19190.4]
  wire  acc_9_io_deq_valid; // @[TensorGemm.scala 156:34:@19190.4]
  wire [31:0] acc_9_io_deq_bits; // @[TensorGemm.scala 156:34:@19190.4]
  wire  acc_10_clock; // @[TensorGemm.scala 156:34:@19193.4]
  wire  acc_10_reset; // @[TensorGemm.scala 156:34:@19193.4]
  wire  acc_10_io_enq_valid; // @[TensorGemm.scala 156:34:@19193.4]
  wire [31:0] acc_10_io_enq_bits; // @[TensorGemm.scala 156:34:@19193.4]
  wire  acc_10_io_deq_valid; // @[TensorGemm.scala 156:34:@19193.4]
  wire [31:0] acc_10_io_deq_bits; // @[TensorGemm.scala 156:34:@19193.4]
  wire  acc_11_clock; // @[TensorGemm.scala 156:34:@19196.4]
  wire  acc_11_reset; // @[TensorGemm.scala 156:34:@19196.4]
  wire  acc_11_io_enq_valid; // @[TensorGemm.scala 156:34:@19196.4]
  wire [31:0] acc_11_io_enq_bits; // @[TensorGemm.scala 156:34:@19196.4]
  wire  acc_11_io_deq_valid; // @[TensorGemm.scala 156:34:@19196.4]
  wire [31:0] acc_11_io_deq_bits; // @[TensorGemm.scala 156:34:@19196.4]
  wire  acc_12_clock; // @[TensorGemm.scala 156:34:@19199.4]
  wire  acc_12_reset; // @[TensorGemm.scala 156:34:@19199.4]
  wire  acc_12_io_enq_valid; // @[TensorGemm.scala 156:34:@19199.4]
  wire [31:0] acc_12_io_enq_bits; // @[TensorGemm.scala 156:34:@19199.4]
  wire  acc_12_io_deq_valid; // @[TensorGemm.scala 156:34:@19199.4]
  wire [31:0] acc_12_io_deq_bits; // @[TensorGemm.scala 156:34:@19199.4]
  wire  acc_13_clock; // @[TensorGemm.scala 156:34:@19202.4]
  wire  acc_13_reset; // @[TensorGemm.scala 156:34:@19202.4]
  wire  acc_13_io_enq_valid; // @[TensorGemm.scala 156:34:@19202.4]
  wire [31:0] acc_13_io_enq_bits; // @[TensorGemm.scala 156:34:@19202.4]
  wire  acc_13_io_deq_valid; // @[TensorGemm.scala 156:34:@19202.4]
  wire [31:0] acc_13_io_deq_bits; // @[TensorGemm.scala 156:34:@19202.4]
  wire  acc_14_clock; // @[TensorGemm.scala 156:34:@19205.4]
  wire  acc_14_reset; // @[TensorGemm.scala 156:34:@19205.4]
  wire  acc_14_io_enq_valid; // @[TensorGemm.scala 156:34:@19205.4]
  wire [31:0] acc_14_io_enq_bits; // @[TensorGemm.scala 156:34:@19205.4]
  wire  acc_14_io_deq_valid; // @[TensorGemm.scala 156:34:@19205.4]
  wire [31:0] acc_14_io_deq_bits; // @[TensorGemm.scala 156:34:@19205.4]
  wire  acc_15_clock; // @[TensorGemm.scala 156:34:@19208.4]
  wire  acc_15_reset; // @[TensorGemm.scala 156:34:@19208.4]
  wire  acc_15_io_enq_valid; // @[TensorGemm.scala 156:34:@19208.4]
  wire [31:0] acc_15_io_enq_bits; // @[TensorGemm.scala 156:34:@19208.4]
  wire  acc_15_io_deq_valid; // @[TensorGemm.scala 156:34:@19208.4]
  wire [31:0] acc_15_io_deq_bits; // @[TensorGemm.scala 156:34:@19208.4]
  wire  _T_6016; // @[TensorGemm.scala 161:46:@19228.4]
  wire  _T_6017; // @[TensorGemm.scala 161:66:@19229.4]
  wire  _T_6018; // @[TensorGemm.scala 161:90:@19230.4]
  wire [31:0] _T_6052; // @[TensorGemm.scala 167:34:@19298.4]
  wire [31:0] _GEN_0; // @[TensorGemm.scala 167:41:@19299.4]
  wire [32:0] _T_6053; // @[TensorGemm.scala 167:41:@19299.4]
  wire [31:0] _T_6054; // @[TensorGemm.scala 167:41:@19300.4]
  wire [31:0] add_0; // @[TensorGemm.scala 167:41:@19301.4]
  wire [31:0] _T_6057; // @[TensorGemm.scala 168:59:@19303.4]
  wire [31:0] _T_6096; // @[TensorGemm.scala 167:34:@19379.4]
  wire [31:0] _GEN_1; // @[TensorGemm.scala 167:41:@19380.4]
  wire [32:0] _T_6097; // @[TensorGemm.scala 167:41:@19380.4]
  wire [31:0] _T_6098; // @[TensorGemm.scala 167:41:@19381.4]
  wire [31:0] add_1; // @[TensorGemm.scala 167:41:@19382.4]
  wire [31:0] _T_6101; // @[TensorGemm.scala 168:59:@19384.4]
  wire [31:0] _T_6140; // @[TensorGemm.scala 167:34:@19460.4]
  wire [31:0] _GEN_2; // @[TensorGemm.scala 167:41:@19461.4]
  wire [32:0] _T_6141; // @[TensorGemm.scala 167:41:@19461.4]
  wire [31:0] _T_6142; // @[TensorGemm.scala 167:41:@19462.4]
  wire [31:0] add_2; // @[TensorGemm.scala 167:41:@19463.4]
  wire [31:0] _T_6145; // @[TensorGemm.scala 168:59:@19465.4]
  wire [31:0] _T_6184; // @[TensorGemm.scala 167:34:@19541.4]
  wire [31:0] _GEN_3; // @[TensorGemm.scala 167:41:@19542.4]
  wire [32:0] _T_6185; // @[TensorGemm.scala 167:41:@19542.4]
  wire [31:0] _T_6186; // @[TensorGemm.scala 167:41:@19543.4]
  wire [31:0] add_3; // @[TensorGemm.scala 167:41:@19544.4]
  wire [31:0] _T_6189; // @[TensorGemm.scala 168:59:@19546.4]
  wire [31:0] _T_6228; // @[TensorGemm.scala 167:34:@19622.4]
  wire [31:0] _GEN_4; // @[TensorGemm.scala 167:41:@19623.4]
  wire [32:0] _T_6229; // @[TensorGemm.scala 167:41:@19623.4]
  wire [31:0] _T_6230; // @[TensorGemm.scala 167:41:@19624.4]
  wire [31:0] add_4; // @[TensorGemm.scala 167:41:@19625.4]
  wire [31:0] _T_6233; // @[TensorGemm.scala 168:59:@19627.4]
  wire [31:0] _T_6272; // @[TensorGemm.scala 167:34:@19703.4]
  wire [31:0] _GEN_5; // @[TensorGemm.scala 167:41:@19704.4]
  wire [32:0] _T_6273; // @[TensorGemm.scala 167:41:@19704.4]
  wire [31:0] _T_6274; // @[TensorGemm.scala 167:41:@19705.4]
  wire [31:0] add_5; // @[TensorGemm.scala 167:41:@19706.4]
  wire [31:0] _T_6277; // @[TensorGemm.scala 168:59:@19708.4]
  wire [31:0] _T_6316; // @[TensorGemm.scala 167:34:@19784.4]
  wire [31:0] _GEN_6; // @[TensorGemm.scala 167:41:@19785.4]
  wire [32:0] _T_6317; // @[TensorGemm.scala 167:41:@19785.4]
  wire [31:0] _T_6318; // @[TensorGemm.scala 167:41:@19786.4]
  wire [31:0] add_6; // @[TensorGemm.scala 167:41:@19787.4]
  wire [31:0] _T_6321; // @[TensorGemm.scala 168:59:@19789.4]
  wire [31:0] _T_6360; // @[TensorGemm.scala 167:34:@19865.4]
  wire [31:0] _GEN_7; // @[TensorGemm.scala 167:41:@19866.4]
  wire [32:0] _T_6361; // @[TensorGemm.scala 167:41:@19866.4]
  wire [31:0] _T_6362; // @[TensorGemm.scala 167:41:@19867.4]
  wire [31:0] add_7; // @[TensorGemm.scala 167:41:@19868.4]
  wire [31:0] _T_6365; // @[TensorGemm.scala 168:59:@19870.4]
  wire [31:0] _T_6404; // @[TensorGemm.scala 167:34:@19946.4]
  wire [31:0] _GEN_8; // @[TensorGemm.scala 167:41:@19947.4]
  wire [32:0] _T_6405; // @[TensorGemm.scala 167:41:@19947.4]
  wire [31:0] _T_6406; // @[TensorGemm.scala 167:41:@19948.4]
  wire [31:0] add_8; // @[TensorGemm.scala 167:41:@19949.4]
  wire [31:0] _T_6409; // @[TensorGemm.scala 168:59:@19951.4]
  wire [31:0] _T_6448; // @[TensorGemm.scala 167:34:@20027.4]
  wire [31:0] _GEN_9; // @[TensorGemm.scala 167:41:@20028.4]
  wire [32:0] _T_6449; // @[TensorGemm.scala 167:41:@20028.4]
  wire [31:0] _T_6450; // @[TensorGemm.scala 167:41:@20029.4]
  wire [31:0] add_9; // @[TensorGemm.scala 167:41:@20030.4]
  wire [31:0] _T_6453; // @[TensorGemm.scala 168:59:@20032.4]
  wire [31:0] _T_6492; // @[TensorGemm.scala 167:34:@20108.4]
  wire [31:0] _GEN_10; // @[TensorGemm.scala 167:41:@20109.4]
  wire [32:0] _T_6493; // @[TensorGemm.scala 167:41:@20109.4]
  wire [31:0] _T_6494; // @[TensorGemm.scala 167:41:@20110.4]
  wire [31:0] add_10; // @[TensorGemm.scala 167:41:@20111.4]
  wire [31:0] _T_6497; // @[TensorGemm.scala 168:59:@20113.4]
  wire [31:0] _T_6536; // @[TensorGemm.scala 167:34:@20189.4]
  wire [31:0] _GEN_11; // @[TensorGemm.scala 167:41:@20190.4]
  wire [32:0] _T_6537; // @[TensorGemm.scala 167:41:@20190.4]
  wire [31:0] _T_6538; // @[TensorGemm.scala 167:41:@20191.4]
  wire [31:0] add_11; // @[TensorGemm.scala 167:41:@20192.4]
  wire [31:0] _T_6541; // @[TensorGemm.scala 168:59:@20194.4]
  wire [31:0] _T_6580; // @[TensorGemm.scala 167:34:@20270.4]
  wire [31:0] _GEN_12; // @[TensorGemm.scala 167:41:@20271.4]
  wire [32:0] _T_6581; // @[TensorGemm.scala 167:41:@20271.4]
  wire [31:0] _T_6582; // @[TensorGemm.scala 167:41:@20272.4]
  wire [31:0] add_12; // @[TensorGemm.scala 167:41:@20273.4]
  wire [31:0] _T_6585; // @[TensorGemm.scala 168:59:@20275.4]
  wire [31:0] _T_6624; // @[TensorGemm.scala 167:34:@20351.4]
  wire [31:0] _GEN_13; // @[TensorGemm.scala 167:41:@20352.4]
  wire [32:0] _T_6625; // @[TensorGemm.scala 167:41:@20352.4]
  wire [31:0] _T_6626; // @[TensorGemm.scala 167:41:@20353.4]
  wire [31:0] add_13; // @[TensorGemm.scala 167:41:@20354.4]
  wire [31:0] _T_6629; // @[TensorGemm.scala 168:59:@20356.4]
  wire [31:0] _T_6668; // @[TensorGemm.scala 167:34:@20432.4]
  wire [31:0] _GEN_14; // @[TensorGemm.scala 167:41:@20433.4]
  wire [32:0] _T_6669; // @[TensorGemm.scala 167:41:@20433.4]
  wire [31:0] _T_6670; // @[TensorGemm.scala 167:41:@20434.4]
  wire [31:0] add_14; // @[TensorGemm.scala 167:41:@20435.4]
  wire [31:0] _T_6673; // @[TensorGemm.scala 168:59:@20437.4]
  wire [31:0] _T_6712; // @[TensorGemm.scala 167:34:@20513.4]
  wire [31:0] _GEN_15; // @[TensorGemm.scala 167:41:@20514.4]
  wire [32:0] _T_6713; // @[TensorGemm.scala 167:41:@20514.4]
  wire [31:0] _T_6714; // @[TensorGemm.scala 167:41:@20515.4]
  wire [31:0] add_15; // @[TensorGemm.scala 167:41:@20516.4]
  wire [31:0] _T_6717; // @[TensorGemm.scala 168:59:@20518.4]
  wire  vld_1; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19389.4]
  wire  vld_0; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19308.4]
  wire  vld_3; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19551.4]
  wire  vld_2; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19470.4]
  wire  vld_5; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19713.4]
  wire  vld_4; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19632.4]
  wire  vld_7; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19875.4]
  wire  vld_6; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19794.4]
  wire [7:0] _T_6726; // @[TensorGemm.scala 172:30:@20530.4]
  wire  vld_9; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20037.4]
  wire  vld_8; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19956.4]
  wire  vld_11; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20199.4]
  wire  vld_10; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20118.4]
  wire  vld_13; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20361.4]
  wire  vld_12; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20280.4]
  wire  vld_15; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20523.4]
  wire  vld_14; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20442.4]
  wire [15:0] _T_6734; // @[TensorGemm.scala 172:30:@20538.4]
  wire [15:0] _T_6735; // @[TensorGemm.scala 172:37:@20539.4]
  wire  _T_6737; // @[TensorGemm.scala 172:37:@20540.4]
  DotProduct dot_0 ( // @[TensorGemm.scala 153:11:@19115.4]
    .clock(dot_0_clock),
    .io_a_0(dot_0_io_a_0),
    .io_a_1(dot_0_io_a_1),
    .io_a_2(dot_0_io_a_2),
    .io_a_3(dot_0_io_a_3),
    .io_a_4(dot_0_io_a_4),
    .io_a_5(dot_0_io_a_5),
    .io_a_6(dot_0_io_a_6),
    .io_a_7(dot_0_io_a_7),
    .io_a_8(dot_0_io_a_8),
    .io_a_9(dot_0_io_a_9),
    .io_a_10(dot_0_io_a_10),
    .io_a_11(dot_0_io_a_11),
    .io_a_12(dot_0_io_a_12),
    .io_a_13(dot_0_io_a_13),
    .io_a_14(dot_0_io_a_14),
    .io_a_15(dot_0_io_a_15),
    .io_b_0(dot_0_io_b_0),
    .io_b_1(dot_0_io_b_1),
    .io_b_2(dot_0_io_b_2),
    .io_b_3(dot_0_io_b_3),
    .io_b_4(dot_0_io_b_4),
    .io_b_5(dot_0_io_b_5),
    .io_b_6(dot_0_io_b_6),
    .io_b_7(dot_0_io_b_7),
    .io_b_8(dot_0_io_b_8),
    .io_b_9(dot_0_io_b_9),
    .io_b_10(dot_0_io_b_10),
    .io_b_11(dot_0_io_b_11),
    .io_b_12(dot_0_io_b_12),
    .io_b_13(dot_0_io_b_13),
    .io_b_14(dot_0_io_b_14),
    .io_b_15(dot_0_io_b_15),
    .io_y(dot_0_io_y)
  );
  DotProduct dot_1 ( // @[TensorGemm.scala 153:11:@19118.4]
    .clock(dot_1_clock),
    .io_a_0(dot_1_io_a_0),
    .io_a_1(dot_1_io_a_1),
    .io_a_2(dot_1_io_a_2),
    .io_a_3(dot_1_io_a_3),
    .io_a_4(dot_1_io_a_4),
    .io_a_5(dot_1_io_a_5),
    .io_a_6(dot_1_io_a_6),
    .io_a_7(dot_1_io_a_7),
    .io_a_8(dot_1_io_a_8),
    .io_a_9(dot_1_io_a_9),
    .io_a_10(dot_1_io_a_10),
    .io_a_11(dot_1_io_a_11),
    .io_a_12(dot_1_io_a_12),
    .io_a_13(dot_1_io_a_13),
    .io_a_14(dot_1_io_a_14),
    .io_a_15(dot_1_io_a_15),
    .io_b_0(dot_1_io_b_0),
    .io_b_1(dot_1_io_b_1),
    .io_b_2(dot_1_io_b_2),
    .io_b_3(dot_1_io_b_3),
    .io_b_4(dot_1_io_b_4),
    .io_b_5(dot_1_io_b_5),
    .io_b_6(dot_1_io_b_6),
    .io_b_7(dot_1_io_b_7),
    .io_b_8(dot_1_io_b_8),
    .io_b_9(dot_1_io_b_9),
    .io_b_10(dot_1_io_b_10),
    .io_b_11(dot_1_io_b_11),
    .io_b_12(dot_1_io_b_12),
    .io_b_13(dot_1_io_b_13),
    .io_b_14(dot_1_io_b_14),
    .io_b_15(dot_1_io_b_15),
    .io_y(dot_1_io_y)
  );
  DotProduct dot_2 ( // @[TensorGemm.scala 153:11:@19121.4]
    .clock(dot_2_clock),
    .io_a_0(dot_2_io_a_0),
    .io_a_1(dot_2_io_a_1),
    .io_a_2(dot_2_io_a_2),
    .io_a_3(dot_2_io_a_3),
    .io_a_4(dot_2_io_a_4),
    .io_a_5(dot_2_io_a_5),
    .io_a_6(dot_2_io_a_6),
    .io_a_7(dot_2_io_a_7),
    .io_a_8(dot_2_io_a_8),
    .io_a_9(dot_2_io_a_9),
    .io_a_10(dot_2_io_a_10),
    .io_a_11(dot_2_io_a_11),
    .io_a_12(dot_2_io_a_12),
    .io_a_13(dot_2_io_a_13),
    .io_a_14(dot_2_io_a_14),
    .io_a_15(dot_2_io_a_15),
    .io_b_0(dot_2_io_b_0),
    .io_b_1(dot_2_io_b_1),
    .io_b_2(dot_2_io_b_2),
    .io_b_3(dot_2_io_b_3),
    .io_b_4(dot_2_io_b_4),
    .io_b_5(dot_2_io_b_5),
    .io_b_6(dot_2_io_b_6),
    .io_b_7(dot_2_io_b_7),
    .io_b_8(dot_2_io_b_8),
    .io_b_9(dot_2_io_b_9),
    .io_b_10(dot_2_io_b_10),
    .io_b_11(dot_2_io_b_11),
    .io_b_12(dot_2_io_b_12),
    .io_b_13(dot_2_io_b_13),
    .io_b_14(dot_2_io_b_14),
    .io_b_15(dot_2_io_b_15),
    .io_y(dot_2_io_y)
  );
  DotProduct dot_3 ( // @[TensorGemm.scala 153:11:@19124.4]
    .clock(dot_3_clock),
    .io_a_0(dot_3_io_a_0),
    .io_a_1(dot_3_io_a_1),
    .io_a_2(dot_3_io_a_2),
    .io_a_3(dot_3_io_a_3),
    .io_a_4(dot_3_io_a_4),
    .io_a_5(dot_3_io_a_5),
    .io_a_6(dot_3_io_a_6),
    .io_a_7(dot_3_io_a_7),
    .io_a_8(dot_3_io_a_8),
    .io_a_9(dot_3_io_a_9),
    .io_a_10(dot_3_io_a_10),
    .io_a_11(dot_3_io_a_11),
    .io_a_12(dot_3_io_a_12),
    .io_a_13(dot_3_io_a_13),
    .io_a_14(dot_3_io_a_14),
    .io_a_15(dot_3_io_a_15),
    .io_b_0(dot_3_io_b_0),
    .io_b_1(dot_3_io_b_1),
    .io_b_2(dot_3_io_b_2),
    .io_b_3(dot_3_io_b_3),
    .io_b_4(dot_3_io_b_4),
    .io_b_5(dot_3_io_b_5),
    .io_b_6(dot_3_io_b_6),
    .io_b_7(dot_3_io_b_7),
    .io_b_8(dot_3_io_b_8),
    .io_b_9(dot_3_io_b_9),
    .io_b_10(dot_3_io_b_10),
    .io_b_11(dot_3_io_b_11),
    .io_b_12(dot_3_io_b_12),
    .io_b_13(dot_3_io_b_13),
    .io_b_14(dot_3_io_b_14),
    .io_b_15(dot_3_io_b_15),
    .io_y(dot_3_io_y)
  );
  DotProduct dot_4 ( // @[TensorGemm.scala 153:11:@19127.4]
    .clock(dot_4_clock),
    .io_a_0(dot_4_io_a_0),
    .io_a_1(dot_4_io_a_1),
    .io_a_2(dot_4_io_a_2),
    .io_a_3(dot_4_io_a_3),
    .io_a_4(dot_4_io_a_4),
    .io_a_5(dot_4_io_a_5),
    .io_a_6(dot_4_io_a_6),
    .io_a_7(dot_4_io_a_7),
    .io_a_8(dot_4_io_a_8),
    .io_a_9(dot_4_io_a_9),
    .io_a_10(dot_4_io_a_10),
    .io_a_11(dot_4_io_a_11),
    .io_a_12(dot_4_io_a_12),
    .io_a_13(dot_4_io_a_13),
    .io_a_14(dot_4_io_a_14),
    .io_a_15(dot_4_io_a_15),
    .io_b_0(dot_4_io_b_0),
    .io_b_1(dot_4_io_b_1),
    .io_b_2(dot_4_io_b_2),
    .io_b_3(dot_4_io_b_3),
    .io_b_4(dot_4_io_b_4),
    .io_b_5(dot_4_io_b_5),
    .io_b_6(dot_4_io_b_6),
    .io_b_7(dot_4_io_b_7),
    .io_b_8(dot_4_io_b_8),
    .io_b_9(dot_4_io_b_9),
    .io_b_10(dot_4_io_b_10),
    .io_b_11(dot_4_io_b_11),
    .io_b_12(dot_4_io_b_12),
    .io_b_13(dot_4_io_b_13),
    .io_b_14(dot_4_io_b_14),
    .io_b_15(dot_4_io_b_15),
    .io_y(dot_4_io_y)
  );
  DotProduct dot_5 ( // @[TensorGemm.scala 153:11:@19130.4]
    .clock(dot_5_clock),
    .io_a_0(dot_5_io_a_0),
    .io_a_1(dot_5_io_a_1),
    .io_a_2(dot_5_io_a_2),
    .io_a_3(dot_5_io_a_3),
    .io_a_4(dot_5_io_a_4),
    .io_a_5(dot_5_io_a_5),
    .io_a_6(dot_5_io_a_6),
    .io_a_7(dot_5_io_a_7),
    .io_a_8(dot_5_io_a_8),
    .io_a_9(dot_5_io_a_9),
    .io_a_10(dot_5_io_a_10),
    .io_a_11(dot_5_io_a_11),
    .io_a_12(dot_5_io_a_12),
    .io_a_13(dot_5_io_a_13),
    .io_a_14(dot_5_io_a_14),
    .io_a_15(dot_5_io_a_15),
    .io_b_0(dot_5_io_b_0),
    .io_b_1(dot_5_io_b_1),
    .io_b_2(dot_5_io_b_2),
    .io_b_3(dot_5_io_b_3),
    .io_b_4(dot_5_io_b_4),
    .io_b_5(dot_5_io_b_5),
    .io_b_6(dot_5_io_b_6),
    .io_b_7(dot_5_io_b_7),
    .io_b_8(dot_5_io_b_8),
    .io_b_9(dot_5_io_b_9),
    .io_b_10(dot_5_io_b_10),
    .io_b_11(dot_5_io_b_11),
    .io_b_12(dot_5_io_b_12),
    .io_b_13(dot_5_io_b_13),
    .io_b_14(dot_5_io_b_14),
    .io_b_15(dot_5_io_b_15),
    .io_y(dot_5_io_y)
  );
  DotProduct dot_6 ( // @[TensorGemm.scala 153:11:@19133.4]
    .clock(dot_6_clock),
    .io_a_0(dot_6_io_a_0),
    .io_a_1(dot_6_io_a_1),
    .io_a_2(dot_6_io_a_2),
    .io_a_3(dot_6_io_a_3),
    .io_a_4(dot_6_io_a_4),
    .io_a_5(dot_6_io_a_5),
    .io_a_6(dot_6_io_a_6),
    .io_a_7(dot_6_io_a_7),
    .io_a_8(dot_6_io_a_8),
    .io_a_9(dot_6_io_a_9),
    .io_a_10(dot_6_io_a_10),
    .io_a_11(dot_6_io_a_11),
    .io_a_12(dot_6_io_a_12),
    .io_a_13(dot_6_io_a_13),
    .io_a_14(dot_6_io_a_14),
    .io_a_15(dot_6_io_a_15),
    .io_b_0(dot_6_io_b_0),
    .io_b_1(dot_6_io_b_1),
    .io_b_2(dot_6_io_b_2),
    .io_b_3(dot_6_io_b_3),
    .io_b_4(dot_6_io_b_4),
    .io_b_5(dot_6_io_b_5),
    .io_b_6(dot_6_io_b_6),
    .io_b_7(dot_6_io_b_7),
    .io_b_8(dot_6_io_b_8),
    .io_b_9(dot_6_io_b_9),
    .io_b_10(dot_6_io_b_10),
    .io_b_11(dot_6_io_b_11),
    .io_b_12(dot_6_io_b_12),
    .io_b_13(dot_6_io_b_13),
    .io_b_14(dot_6_io_b_14),
    .io_b_15(dot_6_io_b_15),
    .io_y(dot_6_io_y)
  );
  DotProduct dot_7 ( // @[TensorGemm.scala 153:11:@19136.4]
    .clock(dot_7_clock),
    .io_a_0(dot_7_io_a_0),
    .io_a_1(dot_7_io_a_1),
    .io_a_2(dot_7_io_a_2),
    .io_a_3(dot_7_io_a_3),
    .io_a_4(dot_7_io_a_4),
    .io_a_5(dot_7_io_a_5),
    .io_a_6(dot_7_io_a_6),
    .io_a_7(dot_7_io_a_7),
    .io_a_8(dot_7_io_a_8),
    .io_a_9(dot_7_io_a_9),
    .io_a_10(dot_7_io_a_10),
    .io_a_11(dot_7_io_a_11),
    .io_a_12(dot_7_io_a_12),
    .io_a_13(dot_7_io_a_13),
    .io_a_14(dot_7_io_a_14),
    .io_a_15(dot_7_io_a_15),
    .io_b_0(dot_7_io_b_0),
    .io_b_1(dot_7_io_b_1),
    .io_b_2(dot_7_io_b_2),
    .io_b_3(dot_7_io_b_3),
    .io_b_4(dot_7_io_b_4),
    .io_b_5(dot_7_io_b_5),
    .io_b_6(dot_7_io_b_6),
    .io_b_7(dot_7_io_b_7),
    .io_b_8(dot_7_io_b_8),
    .io_b_9(dot_7_io_b_9),
    .io_b_10(dot_7_io_b_10),
    .io_b_11(dot_7_io_b_11),
    .io_b_12(dot_7_io_b_12),
    .io_b_13(dot_7_io_b_13),
    .io_b_14(dot_7_io_b_14),
    .io_b_15(dot_7_io_b_15),
    .io_y(dot_7_io_y)
  );
  DotProduct dot_8 ( // @[TensorGemm.scala 153:11:@19139.4]
    .clock(dot_8_clock),
    .io_a_0(dot_8_io_a_0),
    .io_a_1(dot_8_io_a_1),
    .io_a_2(dot_8_io_a_2),
    .io_a_3(dot_8_io_a_3),
    .io_a_4(dot_8_io_a_4),
    .io_a_5(dot_8_io_a_5),
    .io_a_6(dot_8_io_a_6),
    .io_a_7(dot_8_io_a_7),
    .io_a_8(dot_8_io_a_8),
    .io_a_9(dot_8_io_a_9),
    .io_a_10(dot_8_io_a_10),
    .io_a_11(dot_8_io_a_11),
    .io_a_12(dot_8_io_a_12),
    .io_a_13(dot_8_io_a_13),
    .io_a_14(dot_8_io_a_14),
    .io_a_15(dot_8_io_a_15),
    .io_b_0(dot_8_io_b_0),
    .io_b_1(dot_8_io_b_1),
    .io_b_2(dot_8_io_b_2),
    .io_b_3(dot_8_io_b_3),
    .io_b_4(dot_8_io_b_4),
    .io_b_5(dot_8_io_b_5),
    .io_b_6(dot_8_io_b_6),
    .io_b_7(dot_8_io_b_7),
    .io_b_8(dot_8_io_b_8),
    .io_b_9(dot_8_io_b_9),
    .io_b_10(dot_8_io_b_10),
    .io_b_11(dot_8_io_b_11),
    .io_b_12(dot_8_io_b_12),
    .io_b_13(dot_8_io_b_13),
    .io_b_14(dot_8_io_b_14),
    .io_b_15(dot_8_io_b_15),
    .io_y(dot_8_io_y)
  );
  DotProduct dot_9 ( // @[TensorGemm.scala 153:11:@19142.4]
    .clock(dot_9_clock),
    .io_a_0(dot_9_io_a_0),
    .io_a_1(dot_9_io_a_1),
    .io_a_2(dot_9_io_a_2),
    .io_a_3(dot_9_io_a_3),
    .io_a_4(dot_9_io_a_4),
    .io_a_5(dot_9_io_a_5),
    .io_a_6(dot_9_io_a_6),
    .io_a_7(dot_9_io_a_7),
    .io_a_8(dot_9_io_a_8),
    .io_a_9(dot_9_io_a_9),
    .io_a_10(dot_9_io_a_10),
    .io_a_11(dot_9_io_a_11),
    .io_a_12(dot_9_io_a_12),
    .io_a_13(dot_9_io_a_13),
    .io_a_14(dot_9_io_a_14),
    .io_a_15(dot_9_io_a_15),
    .io_b_0(dot_9_io_b_0),
    .io_b_1(dot_9_io_b_1),
    .io_b_2(dot_9_io_b_2),
    .io_b_3(dot_9_io_b_3),
    .io_b_4(dot_9_io_b_4),
    .io_b_5(dot_9_io_b_5),
    .io_b_6(dot_9_io_b_6),
    .io_b_7(dot_9_io_b_7),
    .io_b_8(dot_9_io_b_8),
    .io_b_9(dot_9_io_b_9),
    .io_b_10(dot_9_io_b_10),
    .io_b_11(dot_9_io_b_11),
    .io_b_12(dot_9_io_b_12),
    .io_b_13(dot_9_io_b_13),
    .io_b_14(dot_9_io_b_14),
    .io_b_15(dot_9_io_b_15),
    .io_y(dot_9_io_y)
  );
  DotProduct dot_10 ( // @[TensorGemm.scala 153:11:@19145.4]
    .clock(dot_10_clock),
    .io_a_0(dot_10_io_a_0),
    .io_a_1(dot_10_io_a_1),
    .io_a_2(dot_10_io_a_2),
    .io_a_3(dot_10_io_a_3),
    .io_a_4(dot_10_io_a_4),
    .io_a_5(dot_10_io_a_5),
    .io_a_6(dot_10_io_a_6),
    .io_a_7(dot_10_io_a_7),
    .io_a_8(dot_10_io_a_8),
    .io_a_9(dot_10_io_a_9),
    .io_a_10(dot_10_io_a_10),
    .io_a_11(dot_10_io_a_11),
    .io_a_12(dot_10_io_a_12),
    .io_a_13(dot_10_io_a_13),
    .io_a_14(dot_10_io_a_14),
    .io_a_15(dot_10_io_a_15),
    .io_b_0(dot_10_io_b_0),
    .io_b_1(dot_10_io_b_1),
    .io_b_2(dot_10_io_b_2),
    .io_b_3(dot_10_io_b_3),
    .io_b_4(dot_10_io_b_4),
    .io_b_5(dot_10_io_b_5),
    .io_b_6(dot_10_io_b_6),
    .io_b_7(dot_10_io_b_7),
    .io_b_8(dot_10_io_b_8),
    .io_b_9(dot_10_io_b_9),
    .io_b_10(dot_10_io_b_10),
    .io_b_11(dot_10_io_b_11),
    .io_b_12(dot_10_io_b_12),
    .io_b_13(dot_10_io_b_13),
    .io_b_14(dot_10_io_b_14),
    .io_b_15(dot_10_io_b_15),
    .io_y(dot_10_io_y)
  );
  DotProduct dot_11 ( // @[TensorGemm.scala 153:11:@19148.4]
    .clock(dot_11_clock),
    .io_a_0(dot_11_io_a_0),
    .io_a_1(dot_11_io_a_1),
    .io_a_2(dot_11_io_a_2),
    .io_a_3(dot_11_io_a_3),
    .io_a_4(dot_11_io_a_4),
    .io_a_5(dot_11_io_a_5),
    .io_a_6(dot_11_io_a_6),
    .io_a_7(dot_11_io_a_7),
    .io_a_8(dot_11_io_a_8),
    .io_a_9(dot_11_io_a_9),
    .io_a_10(dot_11_io_a_10),
    .io_a_11(dot_11_io_a_11),
    .io_a_12(dot_11_io_a_12),
    .io_a_13(dot_11_io_a_13),
    .io_a_14(dot_11_io_a_14),
    .io_a_15(dot_11_io_a_15),
    .io_b_0(dot_11_io_b_0),
    .io_b_1(dot_11_io_b_1),
    .io_b_2(dot_11_io_b_2),
    .io_b_3(dot_11_io_b_3),
    .io_b_4(dot_11_io_b_4),
    .io_b_5(dot_11_io_b_5),
    .io_b_6(dot_11_io_b_6),
    .io_b_7(dot_11_io_b_7),
    .io_b_8(dot_11_io_b_8),
    .io_b_9(dot_11_io_b_9),
    .io_b_10(dot_11_io_b_10),
    .io_b_11(dot_11_io_b_11),
    .io_b_12(dot_11_io_b_12),
    .io_b_13(dot_11_io_b_13),
    .io_b_14(dot_11_io_b_14),
    .io_b_15(dot_11_io_b_15),
    .io_y(dot_11_io_y)
  );
  DotProduct dot_12 ( // @[TensorGemm.scala 153:11:@19151.4]
    .clock(dot_12_clock),
    .io_a_0(dot_12_io_a_0),
    .io_a_1(dot_12_io_a_1),
    .io_a_2(dot_12_io_a_2),
    .io_a_3(dot_12_io_a_3),
    .io_a_4(dot_12_io_a_4),
    .io_a_5(dot_12_io_a_5),
    .io_a_6(dot_12_io_a_6),
    .io_a_7(dot_12_io_a_7),
    .io_a_8(dot_12_io_a_8),
    .io_a_9(dot_12_io_a_9),
    .io_a_10(dot_12_io_a_10),
    .io_a_11(dot_12_io_a_11),
    .io_a_12(dot_12_io_a_12),
    .io_a_13(dot_12_io_a_13),
    .io_a_14(dot_12_io_a_14),
    .io_a_15(dot_12_io_a_15),
    .io_b_0(dot_12_io_b_0),
    .io_b_1(dot_12_io_b_1),
    .io_b_2(dot_12_io_b_2),
    .io_b_3(dot_12_io_b_3),
    .io_b_4(dot_12_io_b_4),
    .io_b_5(dot_12_io_b_5),
    .io_b_6(dot_12_io_b_6),
    .io_b_7(dot_12_io_b_7),
    .io_b_8(dot_12_io_b_8),
    .io_b_9(dot_12_io_b_9),
    .io_b_10(dot_12_io_b_10),
    .io_b_11(dot_12_io_b_11),
    .io_b_12(dot_12_io_b_12),
    .io_b_13(dot_12_io_b_13),
    .io_b_14(dot_12_io_b_14),
    .io_b_15(dot_12_io_b_15),
    .io_y(dot_12_io_y)
  );
  DotProduct dot_13 ( // @[TensorGemm.scala 153:11:@19154.4]
    .clock(dot_13_clock),
    .io_a_0(dot_13_io_a_0),
    .io_a_1(dot_13_io_a_1),
    .io_a_2(dot_13_io_a_2),
    .io_a_3(dot_13_io_a_3),
    .io_a_4(dot_13_io_a_4),
    .io_a_5(dot_13_io_a_5),
    .io_a_6(dot_13_io_a_6),
    .io_a_7(dot_13_io_a_7),
    .io_a_8(dot_13_io_a_8),
    .io_a_9(dot_13_io_a_9),
    .io_a_10(dot_13_io_a_10),
    .io_a_11(dot_13_io_a_11),
    .io_a_12(dot_13_io_a_12),
    .io_a_13(dot_13_io_a_13),
    .io_a_14(dot_13_io_a_14),
    .io_a_15(dot_13_io_a_15),
    .io_b_0(dot_13_io_b_0),
    .io_b_1(dot_13_io_b_1),
    .io_b_2(dot_13_io_b_2),
    .io_b_3(dot_13_io_b_3),
    .io_b_4(dot_13_io_b_4),
    .io_b_5(dot_13_io_b_5),
    .io_b_6(dot_13_io_b_6),
    .io_b_7(dot_13_io_b_7),
    .io_b_8(dot_13_io_b_8),
    .io_b_9(dot_13_io_b_9),
    .io_b_10(dot_13_io_b_10),
    .io_b_11(dot_13_io_b_11),
    .io_b_12(dot_13_io_b_12),
    .io_b_13(dot_13_io_b_13),
    .io_b_14(dot_13_io_b_14),
    .io_b_15(dot_13_io_b_15),
    .io_y(dot_13_io_y)
  );
  DotProduct dot_14 ( // @[TensorGemm.scala 153:11:@19157.4]
    .clock(dot_14_clock),
    .io_a_0(dot_14_io_a_0),
    .io_a_1(dot_14_io_a_1),
    .io_a_2(dot_14_io_a_2),
    .io_a_3(dot_14_io_a_3),
    .io_a_4(dot_14_io_a_4),
    .io_a_5(dot_14_io_a_5),
    .io_a_6(dot_14_io_a_6),
    .io_a_7(dot_14_io_a_7),
    .io_a_8(dot_14_io_a_8),
    .io_a_9(dot_14_io_a_9),
    .io_a_10(dot_14_io_a_10),
    .io_a_11(dot_14_io_a_11),
    .io_a_12(dot_14_io_a_12),
    .io_a_13(dot_14_io_a_13),
    .io_a_14(dot_14_io_a_14),
    .io_a_15(dot_14_io_a_15),
    .io_b_0(dot_14_io_b_0),
    .io_b_1(dot_14_io_b_1),
    .io_b_2(dot_14_io_b_2),
    .io_b_3(dot_14_io_b_3),
    .io_b_4(dot_14_io_b_4),
    .io_b_5(dot_14_io_b_5),
    .io_b_6(dot_14_io_b_6),
    .io_b_7(dot_14_io_b_7),
    .io_b_8(dot_14_io_b_8),
    .io_b_9(dot_14_io_b_9),
    .io_b_10(dot_14_io_b_10),
    .io_b_11(dot_14_io_b_11),
    .io_b_12(dot_14_io_b_12),
    .io_b_13(dot_14_io_b_13),
    .io_b_14(dot_14_io_b_14),
    .io_b_15(dot_14_io_b_15),
    .io_y(dot_14_io_y)
  );
  DotProduct dot_15 ( // @[TensorGemm.scala 153:11:@19160.4]
    .clock(dot_15_clock),
    .io_a_0(dot_15_io_a_0),
    .io_a_1(dot_15_io_a_1),
    .io_a_2(dot_15_io_a_2),
    .io_a_3(dot_15_io_a_3),
    .io_a_4(dot_15_io_a_4),
    .io_a_5(dot_15_io_a_5),
    .io_a_6(dot_15_io_a_6),
    .io_a_7(dot_15_io_a_7),
    .io_a_8(dot_15_io_a_8),
    .io_a_9(dot_15_io_a_9),
    .io_a_10(dot_15_io_a_10),
    .io_a_11(dot_15_io_a_11),
    .io_a_12(dot_15_io_a_12),
    .io_a_13(dot_15_io_a_13),
    .io_a_14(dot_15_io_a_14),
    .io_a_15(dot_15_io_a_15),
    .io_b_0(dot_15_io_b_0),
    .io_b_1(dot_15_io_b_1),
    .io_b_2(dot_15_io_b_2),
    .io_b_3(dot_15_io_b_3),
    .io_b_4(dot_15_io_b_4),
    .io_b_5(dot_15_io_b_5),
    .io_b_6(dot_15_io_b_6),
    .io_b_7(dot_15_io_b_7),
    .io_b_8(dot_15_io_b_8),
    .io_b_9(dot_15_io_b_9),
    .io_b_10(dot_15_io_b_10),
    .io_b_11(dot_15_io_b_11),
    .io_b_12(dot_15_io_b_12),
    .io_b_13(dot_15_io_b_13),
    .io_b_14(dot_15_io_b_14),
    .io_b_15(dot_15_io_b_15),
    .io_y(dot_15_io_y)
  );
  Pipe acc_0 ( // @[TensorGemm.scala 156:34:@19163.4]
    .clock(acc_0_clock),
    .reset(acc_0_reset),
    .io_enq_valid(acc_0_io_enq_valid),
    .io_enq_bits(acc_0_io_enq_bits),
    .io_deq_valid(acc_0_io_deq_valid),
    .io_deq_bits(acc_0_io_deq_bits)
  );
  Pipe acc_1 ( // @[TensorGemm.scala 156:34:@19166.4]
    .clock(acc_1_clock),
    .reset(acc_1_reset),
    .io_enq_valid(acc_1_io_enq_valid),
    .io_enq_bits(acc_1_io_enq_bits),
    .io_deq_valid(acc_1_io_deq_valid),
    .io_deq_bits(acc_1_io_deq_bits)
  );
  Pipe acc_2 ( // @[TensorGemm.scala 156:34:@19169.4]
    .clock(acc_2_clock),
    .reset(acc_2_reset),
    .io_enq_valid(acc_2_io_enq_valid),
    .io_enq_bits(acc_2_io_enq_bits),
    .io_deq_valid(acc_2_io_deq_valid),
    .io_deq_bits(acc_2_io_deq_bits)
  );
  Pipe acc_3 ( // @[TensorGemm.scala 156:34:@19172.4]
    .clock(acc_3_clock),
    .reset(acc_3_reset),
    .io_enq_valid(acc_3_io_enq_valid),
    .io_enq_bits(acc_3_io_enq_bits),
    .io_deq_valid(acc_3_io_deq_valid),
    .io_deq_bits(acc_3_io_deq_bits)
  );
  Pipe acc_4 ( // @[TensorGemm.scala 156:34:@19175.4]
    .clock(acc_4_clock),
    .reset(acc_4_reset),
    .io_enq_valid(acc_4_io_enq_valid),
    .io_enq_bits(acc_4_io_enq_bits),
    .io_deq_valid(acc_4_io_deq_valid),
    .io_deq_bits(acc_4_io_deq_bits)
  );
  Pipe acc_5 ( // @[TensorGemm.scala 156:34:@19178.4]
    .clock(acc_5_clock),
    .reset(acc_5_reset),
    .io_enq_valid(acc_5_io_enq_valid),
    .io_enq_bits(acc_5_io_enq_bits),
    .io_deq_valid(acc_5_io_deq_valid),
    .io_deq_bits(acc_5_io_deq_bits)
  );
  Pipe acc_6 ( // @[TensorGemm.scala 156:34:@19181.4]
    .clock(acc_6_clock),
    .reset(acc_6_reset),
    .io_enq_valid(acc_6_io_enq_valid),
    .io_enq_bits(acc_6_io_enq_bits),
    .io_deq_valid(acc_6_io_deq_valid),
    .io_deq_bits(acc_6_io_deq_bits)
  );
  Pipe acc_7 ( // @[TensorGemm.scala 156:34:@19184.4]
    .clock(acc_7_clock),
    .reset(acc_7_reset),
    .io_enq_valid(acc_7_io_enq_valid),
    .io_enq_bits(acc_7_io_enq_bits),
    .io_deq_valid(acc_7_io_deq_valid),
    .io_deq_bits(acc_7_io_deq_bits)
  );
  Pipe acc_8 ( // @[TensorGemm.scala 156:34:@19187.4]
    .clock(acc_8_clock),
    .reset(acc_8_reset),
    .io_enq_valid(acc_8_io_enq_valid),
    .io_enq_bits(acc_8_io_enq_bits),
    .io_deq_valid(acc_8_io_deq_valid),
    .io_deq_bits(acc_8_io_deq_bits)
  );
  Pipe acc_9 ( // @[TensorGemm.scala 156:34:@19190.4]
    .clock(acc_9_clock),
    .reset(acc_9_reset),
    .io_enq_valid(acc_9_io_enq_valid),
    .io_enq_bits(acc_9_io_enq_bits),
    .io_deq_valid(acc_9_io_deq_valid),
    .io_deq_bits(acc_9_io_deq_bits)
  );
  Pipe acc_10 ( // @[TensorGemm.scala 156:34:@19193.4]
    .clock(acc_10_clock),
    .reset(acc_10_reset),
    .io_enq_valid(acc_10_io_enq_valid),
    .io_enq_bits(acc_10_io_enq_bits),
    .io_deq_valid(acc_10_io_deq_valid),
    .io_deq_bits(acc_10_io_deq_bits)
  );
  Pipe acc_11 ( // @[TensorGemm.scala 156:34:@19196.4]
    .clock(acc_11_clock),
    .reset(acc_11_reset),
    .io_enq_valid(acc_11_io_enq_valid),
    .io_enq_bits(acc_11_io_enq_bits),
    .io_deq_valid(acc_11_io_deq_valid),
    .io_deq_bits(acc_11_io_deq_bits)
  );
  Pipe acc_12 ( // @[TensorGemm.scala 156:34:@19199.4]
    .clock(acc_12_clock),
    .reset(acc_12_reset),
    .io_enq_valid(acc_12_io_enq_valid),
    .io_enq_bits(acc_12_io_enq_bits),
    .io_deq_valid(acc_12_io_deq_valid),
    .io_deq_bits(acc_12_io_deq_bits)
  );
  Pipe acc_13 ( // @[TensorGemm.scala 156:34:@19202.4]
    .clock(acc_13_clock),
    .reset(acc_13_reset),
    .io_enq_valid(acc_13_io_enq_valid),
    .io_enq_bits(acc_13_io_enq_bits),
    .io_deq_valid(acc_13_io_deq_valid),
    .io_deq_bits(acc_13_io_deq_bits)
  );
  Pipe acc_14 ( // @[TensorGemm.scala 156:34:@19205.4]
    .clock(acc_14_clock),
    .reset(acc_14_reset),
    .io_enq_valid(acc_14_io_enq_valid),
    .io_enq_bits(acc_14_io_enq_bits),
    .io_deq_valid(acc_14_io_deq_valid),
    .io_deq_bits(acc_14_io_deq_bits)
  );
  Pipe acc_15 ( // @[TensorGemm.scala 156:34:@19208.4]
    .clock(acc_15_clock),
    .reset(acc_15_reset),
    .io_enq_valid(acc_15_io_enq_valid),
    .io_enq_bits(acc_15_io_enq_bits),
    .io_deq_valid(acc_15_io_deq_valid),
    .io_deq_bits(acc_15_io_deq_bits)
  );
  assign _T_6016 = io_inp_data_valid & io_wgt_data_valid; // @[TensorGemm.scala 161:46:@19228.4]
  assign _T_6017 = _T_6016 & io_acc_i_data_valid; // @[TensorGemm.scala 161:66:@19229.4]
  assign _T_6018 = ~ io_reset; // @[TensorGemm.scala 161:90:@19230.4]
  assign _T_6052 = $signed(acc_0_io_deq_bits); // @[TensorGemm.scala 167:34:@19298.4]
  assign _GEN_0 = {{11{dot_0_io_y[20]}},dot_0_io_y}; // @[TensorGemm.scala 167:41:@19299.4]
  assign _T_6053 = $signed(_T_6052) + $signed(_GEN_0); // @[TensorGemm.scala 167:41:@19299.4]
  assign _T_6054 = $signed(_T_6052) + $signed(_GEN_0); // @[TensorGemm.scala 167:41:@19300.4]
  assign add_0 = $signed(_T_6054); // @[TensorGemm.scala 167:41:@19301.4]
  assign _T_6057 = $unsigned(add_0); // @[TensorGemm.scala 168:59:@19303.4]
  assign _T_6096 = $signed(acc_1_io_deq_bits); // @[TensorGemm.scala 167:34:@19379.4]
  assign _GEN_1 = {{11{dot_1_io_y[20]}},dot_1_io_y}; // @[TensorGemm.scala 167:41:@19380.4]
  assign _T_6097 = $signed(_T_6096) + $signed(_GEN_1); // @[TensorGemm.scala 167:41:@19380.4]
  assign _T_6098 = $signed(_T_6096) + $signed(_GEN_1); // @[TensorGemm.scala 167:41:@19381.4]
  assign add_1 = $signed(_T_6098); // @[TensorGemm.scala 167:41:@19382.4]
  assign _T_6101 = $unsigned(add_1); // @[TensorGemm.scala 168:59:@19384.4]
  assign _T_6140 = $signed(acc_2_io_deq_bits); // @[TensorGemm.scala 167:34:@19460.4]
  assign _GEN_2 = {{11{dot_2_io_y[20]}},dot_2_io_y}; // @[TensorGemm.scala 167:41:@19461.4]
  assign _T_6141 = $signed(_T_6140) + $signed(_GEN_2); // @[TensorGemm.scala 167:41:@19461.4]
  assign _T_6142 = $signed(_T_6140) + $signed(_GEN_2); // @[TensorGemm.scala 167:41:@19462.4]
  assign add_2 = $signed(_T_6142); // @[TensorGemm.scala 167:41:@19463.4]
  assign _T_6145 = $unsigned(add_2); // @[TensorGemm.scala 168:59:@19465.4]
  assign _T_6184 = $signed(acc_3_io_deq_bits); // @[TensorGemm.scala 167:34:@19541.4]
  assign _GEN_3 = {{11{dot_3_io_y[20]}},dot_3_io_y}; // @[TensorGemm.scala 167:41:@19542.4]
  assign _T_6185 = $signed(_T_6184) + $signed(_GEN_3); // @[TensorGemm.scala 167:41:@19542.4]
  assign _T_6186 = $signed(_T_6184) + $signed(_GEN_3); // @[TensorGemm.scala 167:41:@19543.4]
  assign add_3 = $signed(_T_6186); // @[TensorGemm.scala 167:41:@19544.4]
  assign _T_6189 = $unsigned(add_3); // @[TensorGemm.scala 168:59:@19546.4]
  assign _T_6228 = $signed(acc_4_io_deq_bits); // @[TensorGemm.scala 167:34:@19622.4]
  assign _GEN_4 = {{11{dot_4_io_y[20]}},dot_4_io_y}; // @[TensorGemm.scala 167:41:@19623.4]
  assign _T_6229 = $signed(_T_6228) + $signed(_GEN_4); // @[TensorGemm.scala 167:41:@19623.4]
  assign _T_6230 = $signed(_T_6228) + $signed(_GEN_4); // @[TensorGemm.scala 167:41:@19624.4]
  assign add_4 = $signed(_T_6230); // @[TensorGemm.scala 167:41:@19625.4]
  assign _T_6233 = $unsigned(add_4); // @[TensorGemm.scala 168:59:@19627.4]
  assign _T_6272 = $signed(acc_5_io_deq_bits); // @[TensorGemm.scala 167:34:@19703.4]
  assign _GEN_5 = {{11{dot_5_io_y[20]}},dot_5_io_y}; // @[TensorGemm.scala 167:41:@19704.4]
  assign _T_6273 = $signed(_T_6272) + $signed(_GEN_5); // @[TensorGemm.scala 167:41:@19704.4]
  assign _T_6274 = $signed(_T_6272) + $signed(_GEN_5); // @[TensorGemm.scala 167:41:@19705.4]
  assign add_5 = $signed(_T_6274); // @[TensorGemm.scala 167:41:@19706.4]
  assign _T_6277 = $unsigned(add_5); // @[TensorGemm.scala 168:59:@19708.4]
  assign _T_6316 = $signed(acc_6_io_deq_bits); // @[TensorGemm.scala 167:34:@19784.4]
  assign _GEN_6 = {{11{dot_6_io_y[20]}},dot_6_io_y}; // @[TensorGemm.scala 167:41:@19785.4]
  assign _T_6317 = $signed(_T_6316) + $signed(_GEN_6); // @[TensorGemm.scala 167:41:@19785.4]
  assign _T_6318 = $signed(_T_6316) + $signed(_GEN_6); // @[TensorGemm.scala 167:41:@19786.4]
  assign add_6 = $signed(_T_6318); // @[TensorGemm.scala 167:41:@19787.4]
  assign _T_6321 = $unsigned(add_6); // @[TensorGemm.scala 168:59:@19789.4]
  assign _T_6360 = $signed(acc_7_io_deq_bits); // @[TensorGemm.scala 167:34:@19865.4]
  assign _GEN_7 = {{11{dot_7_io_y[20]}},dot_7_io_y}; // @[TensorGemm.scala 167:41:@19866.4]
  assign _T_6361 = $signed(_T_6360) + $signed(_GEN_7); // @[TensorGemm.scala 167:41:@19866.4]
  assign _T_6362 = $signed(_T_6360) + $signed(_GEN_7); // @[TensorGemm.scala 167:41:@19867.4]
  assign add_7 = $signed(_T_6362); // @[TensorGemm.scala 167:41:@19868.4]
  assign _T_6365 = $unsigned(add_7); // @[TensorGemm.scala 168:59:@19870.4]
  assign _T_6404 = $signed(acc_8_io_deq_bits); // @[TensorGemm.scala 167:34:@19946.4]
  assign _GEN_8 = {{11{dot_8_io_y[20]}},dot_8_io_y}; // @[TensorGemm.scala 167:41:@19947.4]
  assign _T_6405 = $signed(_T_6404) + $signed(_GEN_8); // @[TensorGemm.scala 167:41:@19947.4]
  assign _T_6406 = $signed(_T_6404) + $signed(_GEN_8); // @[TensorGemm.scala 167:41:@19948.4]
  assign add_8 = $signed(_T_6406); // @[TensorGemm.scala 167:41:@19949.4]
  assign _T_6409 = $unsigned(add_8); // @[TensorGemm.scala 168:59:@19951.4]
  assign _T_6448 = $signed(acc_9_io_deq_bits); // @[TensorGemm.scala 167:34:@20027.4]
  assign _GEN_9 = {{11{dot_9_io_y[20]}},dot_9_io_y}; // @[TensorGemm.scala 167:41:@20028.4]
  assign _T_6449 = $signed(_T_6448) + $signed(_GEN_9); // @[TensorGemm.scala 167:41:@20028.4]
  assign _T_6450 = $signed(_T_6448) + $signed(_GEN_9); // @[TensorGemm.scala 167:41:@20029.4]
  assign add_9 = $signed(_T_6450); // @[TensorGemm.scala 167:41:@20030.4]
  assign _T_6453 = $unsigned(add_9); // @[TensorGemm.scala 168:59:@20032.4]
  assign _T_6492 = $signed(acc_10_io_deq_bits); // @[TensorGemm.scala 167:34:@20108.4]
  assign _GEN_10 = {{11{dot_10_io_y[20]}},dot_10_io_y}; // @[TensorGemm.scala 167:41:@20109.4]
  assign _T_6493 = $signed(_T_6492) + $signed(_GEN_10); // @[TensorGemm.scala 167:41:@20109.4]
  assign _T_6494 = $signed(_T_6492) + $signed(_GEN_10); // @[TensorGemm.scala 167:41:@20110.4]
  assign add_10 = $signed(_T_6494); // @[TensorGemm.scala 167:41:@20111.4]
  assign _T_6497 = $unsigned(add_10); // @[TensorGemm.scala 168:59:@20113.4]
  assign _T_6536 = $signed(acc_11_io_deq_bits); // @[TensorGemm.scala 167:34:@20189.4]
  assign _GEN_11 = {{11{dot_11_io_y[20]}},dot_11_io_y}; // @[TensorGemm.scala 167:41:@20190.4]
  assign _T_6537 = $signed(_T_6536) + $signed(_GEN_11); // @[TensorGemm.scala 167:41:@20190.4]
  assign _T_6538 = $signed(_T_6536) + $signed(_GEN_11); // @[TensorGemm.scala 167:41:@20191.4]
  assign add_11 = $signed(_T_6538); // @[TensorGemm.scala 167:41:@20192.4]
  assign _T_6541 = $unsigned(add_11); // @[TensorGemm.scala 168:59:@20194.4]
  assign _T_6580 = $signed(acc_12_io_deq_bits); // @[TensorGemm.scala 167:34:@20270.4]
  assign _GEN_12 = {{11{dot_12_io_y[20]}},dot_12_io_y}; // @[TensorGemm.scala 167:41:@20271.4]
  assign _T_6581 = $signed(_T_6580) + $signed(_GEN_12); // @[TensorGemm.scala 167:41:@20271.4]
  assign _T_6582 = $signed(_T_6580) + $signed(_GEN_12); // @[TensorGemm.scala 167:41:@20272.4]
  assign add_12 = $signed(_T_6582); // @[TensorGemm.scala 167:41:@20273.4]
  assign _T_6585 = $unsigned(add_12); // @[TensorGemm.scala 168:59:@20275.4]
  assign _T_6624 = $signed(acc_13_io_deq_bits); // @[TensorGemm.scala 167:34:@20351.4]
  assign _GEN_13 = {{11{dot_13_io_y[20]}},dot_13_io_y}; // @[TensorGemm.scala 167:41:@20352.4]
  assign _T_6625 = $signed(_T_6624) + $signed(_GEN_13); // @[TensorGemm.scala 167:41:@20352.4]
  assign _T_6626 = $signed(_T_6624) + $signed(_GEN_13); // @[TensorGemm.scala 167:41:@20353.4]
  assign add_13 = $signed(_T_6626); // @[TensorGemm.scala 167:41:@20354.4]
  assign _T_6629 = $unsigned(add_13); // @[TensorGemm.scala 168:59:@20356.4]
  assign _T_6668 = $signed(acc_14_io_deq_bits); // @[TensorGemm.scala 167:34:@20432.4]
  assign _GEN_14 = {{11{dot_14_io_y[20]}},dot_14_io_y}; // @[TensorGemm.scala 167:41:@20433.4]
  assign _T_6669 = $signed(_T_6668) + $signed(_GEN_14); // @[TensorGemm.scala 167:41:@20433.4]
  assign _T_6670 = $signed(_T_6668) + $signed(_GEN_14); // @[TensorGemm.scala 167:41:@20434.4]
  assign add_14 = $signed(_T_6670); // @[TensorGemm.scala 167:41:@20435.4]
  assign _T_6673 = $unsigned(add_14); // @[TensorGemm.scala 168:59:@20437.4]
  assign _T_6712 = $signed(acc_15_io_deq_bits); // @[TensorGemm.scala 167:34:@20513.4]
  assign _GEN_15 = {{11{dot_15_io_y[20]}},dot_15_io_y}; // @[TensorGemm.scala 167:41:@20514.4]
  assign _T_6713 = $signed(_T_6712) + $signed(_GEN_15); // @[TensorGemm.scala 167:41:@20514.4]
  assign _T_6714 = $signed(_T_6712) + $signed(_GEN_15); // @[TensorGemm.scala 167:41:@20515.4]
  assign add_15 = $signed(_T_6714); // @[TensorGemm.scala 167:41:@20516.4]
  assign _T_6717 = $unsigned(add_15); // @[TensorGemm.scala 168:59:@20518.4]
  assign vld_1 = acc_1_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19389.4]
  assign vld_0 = acc_0_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19308.4]
  assign vld_3 = acc_3_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19551.4]
  assign vld_2 = acc_2_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19470.4]
  assign vld_5 = acc_5_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19713.4]
  assign vld_4 = acc_4_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19632.4]
  assign vld_7 = acc_7_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19875.4]
  assign vld_6 = acc_6_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19794.4]
  assign _T_6726 = {vld_7,vld_6,vld_5,vld_4,vld_3,vld_2,vld_1,vld_0}; // @[TensorGemm.scala 172:30:@20530.4]
  assign vld_9 = acc_9_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20037.4]
  assign vld_8 = acc_8_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@19956.4]
  assign vld_11 = acc_11_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20199.4]
  assign vld_10 = acc_10_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20118.4]
  assign vld_13 = acc_13_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20361.4]
  assign vld_12 = acc_12_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20280.4]
  assign vld_15 = acc_15_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20523.4]
  assign vld_14 = acc_14_io_deq_valid; // @[TensorGemm.scala 158:17:@19227.4 TensorGemm.scala 170:12:@20442.4]
  assign _T_6734 = {vld_15,vld_14,vld_13,vld_12,vld_11,vld_10,vld_9,vld_8,_T_6726}; // @[TensorGemm.scala 172:30:@20538.4]
  assign _T_6735 = ~ _T_6734; // @[TensorGemm.scala 172:37:@20539.4]
  assign _T_6737 = _T_6735 == 16'h0; // @[TensorGemm.scala 172:37:@20540.4]
  assign io_acc_o_data_valid = _T_6737 | io_reset; // @[TensorGemm.scala 172:23:@20542.4]
  assign io_acc_o_data_bits_0_0 = io_reset ? 32'h0 : _T_6057; // @[TensorGemm.scala 168:30:@19305.4]
  assign io_acc_o_data_bits_0_1 = io_reset ? 32'h0 : _T_6101; // @[TensorGemm.scala 168:30:@19386.4]
  assign io_acc_o_data_bits_0_2 = io_reset ? 32'h0 : _T_6145; // @[TensorGemm.scala 168:30:@19467.4]
  assign io_acc_o_data_bits_0_3 = io_reset ? 32'h0 : _T_6189; // @[TensorGemm.scala 168:30:@19548.4]
  assign io_acc_o_data_bits_0_4 = io_reset ? 32'h0 : _T_6233; // @[TensorGemm.scala 168:30:@19629.4]
  assign io_acc_o_data_bits_0_5 = io_reset ? 32'h0 : _T_6277; // @[TensorGemm.scala 168:30:@19710.4]
  assign io_acc_o_data_bits_0_6 = io_reset ? 32'h0 : _T_6321; // @[TensorGemm.scala 168:30:@19791.4]
  assign io_acc_o_data_bits_0_7 = io_reset ? 32'h0 : _T_6365; // @[TensorGemm.scala 168:30:@19872.4]
  assign io_acc_o_data_bits_0_8 = io_reset ? 32'h0 : _T_6409; // @[TensorGemm.scala 168:30:@19953.4]
  assign io_acc_o_data_bits_0_9 = io_reset ? 32'h0 : _T_6453; // @[TensorGemm.scala 168:30:@20034.4]
  assign io_acc_o_data_bits_0_10 = io_reset ? 32'h0 : _T_6497; // @[TensorGemm.scala 168:30:@20115.4]
  assign io_acc_o_data_bits_0_11 = io_reset ? 32'h0 : _T_6541; // @[TensorGemm.scala 168:30:@20196.4]
  assign io_acc_o_data_bits_0_12 = io_reset ? 32'h0 : _T_6585; // @[TensorGemm.scala 168:30:@20277.4]
  assign io_acc_o_data_bits_0_13 = io_reset ? 32'h0 : _T_6629; // @[TensorGemm.scala 168:30:@20358.4]
  assign io_acc_o_data_bits_0_14 = io_reset ? 32'h0 : _T_6673; // @[TensorGemm.scala 168:30:@20439.4]
  assign io_acc_o_data_bits_0_15 = io_reset ? 32'h0 : _T_6717; // @[TensorGemm.scala 168:30:@20520.4]
  assign io_out_data_valid = _T_6735 == 16'h0; // @[TensorGemm.scala 173:21:@20560.4]
  assign io_out_data_bits_0_0 = _T_6057[7:0]; // @[TensorGemm.scala 169:28:@19307.4]
  assign io_out_data_bits_0_1 = _T_6101[7:0]; // @[TensorGemm.scala 169:28:@19388.4]
  assign io_out_data_bits_0_2 = _T_6145[7:0]; // @[TensorGemm.scala 169:28:@19469.4]
  assign io_out_data_bits_0_3 = _T_6189[7:0]; // @[TensorGemm.scala 169:28:@19550.4]
  assign io_out_data_bits_0_4 = _T_6233[7:0]; // @[TensorGemm.scala 169:28:@19631.4]
  assign io_out_data_bits_0_5 = _T_6277[7:0]; // @[TensorGemm.scala 169:28:@19712.4]
  assign io_out_data_bits_0_6 = _T_6321[7:0]; // @[TensorGemm.scala 169:28:@19793.4]
  assign io_out_data_bits_0_7 = _T_6365[7:0]; // @[TensorGemm.scala 169:28:@19874.4]
  assign io_out_data_bits_0_8 = _T_6409[7:0]; // @[TensorGemm.scala 169:28:@19955.4]
  assign io_out_data_bits_0_9 = _T_6453[7:0]; // @[TensorGemm.scala 169:28:@20036.4]
  assign io_out_data_bits_0_10 = _T_6497[7:0]; // @[TensorGemm.scala 169:28:@20117.4]
  assign io_out_data_bits_0_11 = _T_6541[7:0]; // @[TensorGemm.scala 169:28:@20198.4]
  assign io_out_data_bits_0_12 = _T_6585[7:0]; // @[TensorGemm.scala 169:28:@20279.4]
  assign io_out_data_bits_0_13 = _T_6629[7:0]; // @[TensorGemm.scala 169:28:@20360.4]
  assign io_out_data_bits_0_14 = _T_6673[7:0]; // @[TensorGemm.scala 169:28:@20441.4]
  assign io_out_data_bits_0_15 = _T_6717[7:0]; // @[TensorGemm.scala 169:28:@20522.4]
  assign dot_0_clock = clock; // @[:@19116.4]
  assign dot_0_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19235.4]
  assign dot_0_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19239.4]
  assign dot_0_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19243.4]
  assign dot_0_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19247.4]
  assign dot_0_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19251.4]
  assign dot_0_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19255.4]
  assign dot_0_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19259.4]
  assign dot_0_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19263.4]
  assign dot_0_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19267.4]
  assign dot_0_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19271.4]
  assign dot_0_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19275.4]
  assign dot_0_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19279.4]
  assign dot_0_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19283.4]
  assign dot_0_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19287.4]
  assign dot_0_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19291.4]
  assign dot_0_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19295.4]
  assign dot_0_io_b_0 = $signed(io_wgt_data_bits_0_0); // @[TensorGemm.scala 165:22:@19237.4]
  assign dot_0_io_b_1 = $signed(io_wgt_data_bits_0_1); // @[TensorGemm.scala 165:22:@19241.4]
  assign dot_0_io_b_2 = $signed(io_wgt_data_bits_0_2); // @[TensorGemm.scala 165:22:@19245.4]
  assign dot_0_io_b_3 = $signed(io_wgt_data_bits_0_3); // @[TensorGemm.scala 165:22:@19249.4]
  assign dot_0_io_b_4 = $signed(io_wgt_data_bits_0_4); // @[TensorGemm.scala 165:22:@19253.4]
  assign dot_0_io_b_5 = $signed(io_wgt_data_bits_0_5); // @[TensorGemm.scala 165:22:@19257.4]
  assign dot_0_io_b_6 = $signed(io_wgt_data_bits_0_6); // @[TensorGemm.scala 165:22:@19261.4]
  assign dot_0_io_b_7 = $signed(io_wgt_data_bits_0_7); // @[TensorGemm.scala 165:22:@19265.4]
  assign dot_0_io_b_8 = $signed(io_wgt_data_bits_0_8); // @[TensorGemm.scala 165:22:@19269.4]
  assign dot_0_io_b_9 = $signed(io_wgt_data_bits_0_9); // @[TensorGemm.scala 165:22:@19273.4]
  assign dot_0_io_b_10 = $signed(io_wgt_data_bits_0_10); // @[TensorGemm.scala 165:22:@19277.4]
  assign dot_0_io_b_11 = $signed(io_wgt_data_bits_0_11); // @[TensorGemm.scala 165:22:@19281.4]
  assign dot_0_io_b_12 = $signed(io_wgt_data_bits_0_12); // @[TensorGemm.scala 165:22:@19285.4]
  assign dot_0_io_b_13 = $signed(io_wgt_data_bits_0_13); // @[TensorGemm.scala 165:22:@19289.4]
  assign dot_0_io_b_14 = $signed(io_wgt_data_bits_0_14); // @[TensorGemm.scala 165:22:@19293.4]
  assign dot_0_io_b_15 = $signed(io_wgt_data_bits_0_15); // @[TensorGemm.scala 165:22:@19297.4]
  assign dot_1_clock = clock; // @[:@19119.4]
  assign dot_1_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19316.4]
  assign dot_1_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19320.4]
  assign dot_1_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19324.4]
  assign dot_1_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19328.4]
  assign dot_1_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19332.4]
  assign dot_1_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19336.4]
  assign dot_1_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19340.4]
  assign dot_1_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19344.4]
  assign dot_1_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19348.4]
  assign dot_1_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19352.4]
  assign dot_1_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19356.4]
  assign dot_1_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19360.4]
  assign dot_1_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19364.4]
  assign dot_1_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19368.4]
  assign dot_1_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19372.4]
  assign dot_1_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19376.4]
  assign dot_1_io_b_0 = $signed(io_wgt_data_bits_1_0); // @[TensorGemm.scala 165:22:@19318.4]
  assign dot_1_io_b_1 = $signed(io_wgt_data_bits_1_1); // @[TensorGemm.scala 165:22:@19322.4]
  assign dot_1_io_b_2 = $signed(io_wgt_data_bits_1_2); // @[TensorGemm.scala 165:22:@19326.4]
  assign dot_1_io_b_3 = $signed(io_wgt_data_bits_1_3); // @[TensorGemm.scala 165:22:@19330.4]
  assign dot_1_io_b_4 = $signed(io_wgt_data_bits_1_4); // @[TensorGemm.scala 165:22:@19334.4]
  assign dot_1_io_b_5 = $signed(io_wgt_data_bits_1_5); // @[TensorGemm.scala 165:22:@19338.4]
  assign dot_1_io_b_6 = $signed(io_wgt_data_bits_1_6); // @[TensorGemm.scala 165:22:@19342.4]
  assign dot_1_io_b_7 = $signed(io_wgt_data_bits_1_7); // @[TensorGemm.scala 165:22:@19346.4]
  assign dot_1_io_b_8 = $signed(io_wgt_data_bits_1_8); // @[TensorGemm.scala 165:22:@19350.4]
  assign dot_1_io_b_9 = $signed(io_wgt_data_bits_1_9); // @[TensorGemm.scala 165:22:@19354.4]
  assign dot_1_io_b_10 = $signed(io_wgt_data_bits_1_10); // @[TensorGemm.scala 165:22:@19358.4]
  assign dot_1_io_b_11 = $signed(io_wgt_data_bits_1_11); // @[TensorGemm.scala 165:22:@19362.4]
  assign dot_1_io_b_12 = $signed(io_wgt_data_bits_1_12); // @[TensorGemm.scala 165:22:@19366.4]
  assign dot_1_io_b_13 = $signed(io_wgt_data_bits_1_13); // @[TensorGemm.scala 165:22:@19370.4]
  assign dot_1_io_b_14 = $signed(io_wgt_data_bits_1_14); // @[TensorGemm.scala 165:22:@19374.4]
  assign dot_1_io_b_15 = $signed(io_wgt_data_bits_1_15); // @[TensorGemm.scala 165:22:@19378.4]
  assign dot_2_clock = clock; // @[:@19122.4]
  assign dot_2_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19397.4]
  assign dot_2_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19401.4]
  assign dot_2_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19405.4]
  assign dot_2_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19409.4]
  assign dot_2_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19413.4]
  assign dot_2_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19417.4]
  assign dot_2_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19421.4]
  assign dot_2_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19425.4]
  assign dot_2_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19429.4]
  assign dot_2_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19433.4]
  assign dot_2_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19437.4]
  assign dot_2_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19441.4]
  assign dot_2_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19445.4]
  assign dot_2_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19449.4]
  assign dot_2_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19453.4]
  assign dot_2_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19457.4]
  assign dot_2_io_b_0 = $signed(io_wgt_data_bits_2_0); // @[TensorGemm.scala 165:22:@19399.4]
  assign dot_2_io_b_1 = $signed(io_wgt_data_bits_2_1); // @[TensorGemm.scala 165:22:@19403.4]
  assign dot_2_io_b_2 = $signed(io_wgt_data_bits_2_2); // @[TensorGemm.scala 165:22:@19407.4]
  assign dot_2_io_b_3 = $signed(io_wgt_data_bits_2_3); // @[TensorGemm.scala 165:22:@19411.4]
  assign dot_2_io_b_4 = $signed(io_wgt_data_bits_2_4); // @[TensorGemm.scala 165:22:@19415.4]
  assign dot_2_io_b_5 = $signed(io_wgt_data_bits_2_5); // @[TensorGemm.scala 165:22:@19419.4]
  assign dot_2_io_b_6 = $signed(io_wgt_data_bits_2_6); // @[TensorGemm.scala 165:22:@19423.4]
  assign dot_2_io_b_7 = $signed(io_wgt_data_bits_2_7); // @[TensorGemm.scala 165:22:@19427.4]
  assign dot_2_io_b_8 = $signed(io_wgt_data_bits_2_8); // @[TensorGemm.scala 165:22:@19431.4]
  assign dot_2_io_b_9 = $signed(io_wgt_data_bits_2_9); // @[TensorGemm.scala 165:22:@19435.4]
  assign dot_2_io_b_10 = $signed(io_wgt_data_bits_2_10); // @[TensorGemm.scala 165:22:@19439.4]
  assign dot_2_io_b_11 = $signed(io_wgt_data_bits_2_11); // @[TensorGemm.scala 165:22:@19443.4]
  assign dot_2_io_b_12 = $signed(io_wgt_data_bits_2_12); // @[TensorGemm.scala 165:22:@19447.4]
  assign dot_2_io_b_13 = $signed(io_wgt_data_bits_2_13); // @[TensorGemm.scala 165:22:@19451.4]
  assign dot_2_io_b_14 = $signed(io_wgt_data_bits_2_14); // @[TensorGemm.scala 165:22:@19455.4]
  assign dot_2_io_b_15 = $signed(io_wgt_data_bits_2_15); // @[TensorGemm.scala 165:22:@19459.4]
  assign dot_3_clock = clock; // @[:@19125.4]
  assign dot_3_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19478.4]
  assign dot_3_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19482.4]
  assign dot_3_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19486.4]
  assign dot_3_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19490.4]
  assign dot_3_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19494.4]
  assign dot_3_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19498.4]
  assign dot_3_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19502.4]
  assign dot_3_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19506.4]
  assign dot_3_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19510.4]
  assign dot_3_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19514.4]
  assign dot_3_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19518.4]
  assign dot_3_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19522.4]
  assign dot_3_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19526.4]
  assign dot_3_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19530.4]
  assign dot_3_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19534.4]
  assign dot_3_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19538.4]
  assign dot_3_io_b_0 = $signed(io_wgt_data_bits_3_0); // @[TensorGemm.scala 165:22:@19480.4]
  assign dot_3_io_b_1 = $signed(io_wgt_data_bits_3_1); // @[TensorGemm.scala 165:22:@19484.4]
  assign dot_3_io_b_2 = $signed(io_wgt_data_bits_3_2); // @[TensorGemm.scala 165:22:@19488.4]
  assign dot_3_io_b_3 = $signed(io_wgt_data_bits_3_3); // @[TensorGemm.scala 165:22:@19492.4]
  assign dot_3_io_b_4 = $signed(io_wgt_data_bits_3_4); // @[TensorGemm.scala 165:22:@19496.4]
  assign dot_3_io_b_5 = $signed(io_wgt_data_bits_3_5); // @[TensorGemm.scala 165:22:@19500.4]
  assign dot_3_io_b_6 = $signed(io_wgt_data_bits_3_6); // @[TensorGemm.scala 165:22:@19504.4]
  assign dot_3_io_b_7 = $signed(io_wgt_data_bits_3_7); // @[TensorGemm.scala 165:22:@19508.4]
  assign dot_3_io_b_8 = $signed(io_wgt_data_bits_3_8); // @[TensorGemm.scala 165:22:@19512.4]
  assign dot_3_io_b_9 = $signed(io_wgt_data_bits_3_9); // @[TensorGemm.scala 165:22:@19516.4]
  assign dot_3_io_b_10 = $signed(io_wgt_data_bits_3_10); // @[TensorGemm.scala 165:22:@19520.4]
  assign dot_3_io_b_11 = $signed(io_wgt_data_bits_3_11); // @[TensorGemm.scala 165:22:@19524.4]
  assign dot_3_io_b_12 = $signed(io_wgt_data_bits_3_12); // @[TensorGemm.scala 165:22:@19528.4]
  assign dot_3_io_b_13 = $signed(io_wgt_data_bits_3_13); // @[TensorGemm.scala 165:22:@19532.4]
  assign dot_3_io_b_14 = $signed(io_wgt_data_bits_3_14); // @[TensorGemm.scala 165:22:@19536.4]
  assign dot_3_io_b_15 = $signed(io_wgt_data_bits_3_15); // @[TensorGemm.scala 165:22:@19540.4]
  assign dot_4_clock = clock; // @[:@19128.4]
  assign dot_4_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19559.4]
  assign dot_4_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19563.4]
  assign dot_4_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19567.4]
  assign dot_4_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19571.4]
  assign dot_4_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19575.4]
  assign dot_4_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19579.4]
  assign dot_4_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19583.4]
  assign dot_4_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19587.4]
  assign dot_4_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19591.4]
  assign dot_4_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19595.4]
  assign dot_4_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19599.4]
  assign dot_4_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19603.4]
  assign dot_4_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19607.4]
  assign dot_4_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19611.4]
  assign dot_4_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19615.4]
  assign dot_4_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19619.4]
  assign dot_4_io_b_0 = $signed(io_wgt_data_bits_4_0); // @[TensorGemm.scala 165:22:@19561.4]
  assign dot_4_io_b_1 = $signed(io_wgt_data_bits_4_1); // @[TensorGemm.scala 165:22:@19565.4]
  assign dot_4_io_b_2 = $signed(io_wgt_data_bits_4_2); // @[TensorGemm.scala 165:22:@19569.4]
  assign dot_4_io_b_3 = $signed(io_wgt_data_bits_4_3); // @[TensorGemm.scala 165:22:@19573.4]
  assign dot_4_io_b_4 = $signed(io_wgt_data_bits_4_4); // @[TensorGemm.scala 165:22:@19577.4]
  assign dot_4_io_b_5 = $signed(io_wgt_data_bits_4_5); // @[TensorGemm.scala 165:22:@19581.4]
  assign dot_4_io_b_6 = $signed(io_wgt_data_bits_4_6); // @[TensorGemm.scala 165:22:@19585.4]
  assign dot_4_io_b_7 = $signed(io_wgt_data_bits_4_7); // @[TensorGemm.scala 165:22:@19589.4]
  assign dot_4_io_b_8 = $signed(io_wgt_data_bits_4_8); // @[TensorGemm.scala 165:22:@19593.4]
  assign dot_4_io_b_9 = $signed(io_wgt_data_bits_4_9); // @[TensorGemm.scala 165:22:@19597.4]
  assign dot_4_io_b_10 = $signed(io_wgt_data_bits_4_10); // @[TensorGemm.scala 165:22:@19601.4]
  assign dot_4_io_b_11 = $signed(io_wgt_data_bits_4_11); // @[TensorGemm.scala 165:22:@19605.4]
  assign dot_4_io_b_12 = $signed(io_wgt_data_bits_4_12); // @[TensorGemm.scala 165:22:@19609.4]
  assign dot_4_io_b_13 = $signed(io_wgt_data_bits_4_13); // @[TensorGemm.scala 165:22:@19613.4]
  assign dot_4_io_b_14 = $signed(io_wgt_data_bits_4_14); // @[TensorGemm.scala 165:22:@19617.4]
  assign dot_4_io_b_15 = $signed(io_wgt_data_bits_4_15); // @[TensorGemm.scala 165:22:@19621.4]
  assign dot_5_clock = clock; // @[:@19131.4]
  assign dot_5_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19640.4]
  assign dot_5_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19644.4]
  assign dot_5_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19648.4]
  assign dot_5_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19652.4]
  assign dot_5_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19656.4]
  assign dot_5_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19660.4]
  assign dot_5_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19664.4]
  assign dot_5_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19668.4]
  assign dot_5_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19672.4]
  assign dot_5_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19676.4]
  assign dot_5_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19680.4]
  assign dot_5_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19684.4]
  assign dot_5_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19688.4]
  assign dot_5_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19692.4]
  assign dot_5_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19696.4]
  assign dot_5_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19700.4]
  assign dot_5_io_b_0 = $signed(io_wgt_data_bits_5_0); // @[TensorGemm.scala 165:22:@19642.4]
  assign dot_5_io_b_1 = $signed(io_wgt_data_bits_5_1); // @[TensorGemm.scala 165:22:@19646.4]
  assign dot_5_io_b_2 = $signed(io_wgt_data_bits_5_2); // @[TensorGemm.scala 165:22:@19650.4]
  assign dot_5_io_b_3 = $signed(io_wgt_data_bits_5_3); // @[TensorGemm.scala 165:22:@19654.4]
  assign dot_5_io_b_4 = $signed(io_wgt_data_bits_5_4); // @[TensorGemm.scala 165:22:@19658.4]
  assign dot_5_io_b_5 = $signed(io_wgt_data_bits_5_5); // @[TensorGemm.scala 165:22:@19662.4]
  assign dot_5_io_b_6 = $signed(io_wgt_data_bits_5_6); // @[TensorGemm.scala 165:22:@19666.4]
  assign dot_5_io_b_7 = $signed(io_wgt_data_bits_5_7); // @[TensorGemm.scala 165:22:@19670.4]
  assign dot_5_io_b_8 = $signed(io_wgt_data_bits_5_8); // @[TensorGemm.scala 165:22:@19674.4]
  assign dot_5_io_b_9 = $signed(io_wgt_data_bits_5_9); // @[TensorGemm.scala 165:22:@19678.4]
  assign dot_5_io_b_10 = $signed(io_wgt_data_bits_5_10); // @[TensorGemm.scala 165:22:@19682.4]
  assign dot_5_io_b_11 = $signed(io_wgt_data_bits_5_11); // @[TensorGemm.scala 165:22:@19686.4]
  assign dot_5_io_b_12 = $signed(io_wgt_data_bits_5_12); // @[TensorGemm.scala 165:22:@19690.4]
  assign dot_5_io_b_13 = $signed(io_wgt_data_bits_5_13); // @[TensorGemm.scala 165:22:@19694.4]
  assign dot_5_io_b_14 = $signed(io_wgt_data_bits_5_14); // @[TensorGemm.scala 165:22:@19698.4]
  assign dot_5_io_b_15 = $signed(io_wgt_data_bits_5_15); // @[TensorGemm.scala 165:22:@19702.4]
  assign dot_6_clock = clock; // @[:@19134.4]
  assign dot_6_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19721.4]
  assign dot_6_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19725.4]
  assign dot_6_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19729.4]
  assign dot_6_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19733.4]
  assign dot_6_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19737.4]
  assign dot_6_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19741.4]
  assign dot_6_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19745.4]
  assign dot_6_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19749.4]
  assign dot_6_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19753.4]
  assign dot_6_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19757.4]
  assign dot_6_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19761.4]
  assign dot_6_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19765.4]
  assign dot_6_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19769.4]
  assign dot_6_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19773.4]
  assign dot_6_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19777.4]
  assign dot_6_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19781.4]
  assign dot_6_io_b_0 = $signed(io_wgt_data_bits_6_0); // @[TensorGemm.scala 165:22:@19723.4]
  assign dot_6_io_b_1 = $signed(io_wgt_data_bits_6_1); // @[TensorGemm.scala 165:22:@19727.4]
  assign dot_6_io_b_2 = $signed(io_wgt_data_bits_6_2); // @[TensorGemm.scala 165:22:@19731.4]
  assign dot_6_io_b_3 = $signed(io_wgt_data_bits_6_3); // @[TensorGemm.scala 165:22:@19735.4]
  assign dot_6_io_b_4 = $signed(io_wgt_data_bits_6_4); // @[TensorGemm.scala 165:22:@19739.4]
  assign dot_6_io_b_5 = $signed(io_wgt_data_bits_6_5); // @[TensorGemm.scala 165:22:@19743.4]
  assign dot_6_io_b_6 = $signed(io_wgt_data_bits_6_6); // @[TensorGemm.scala 165:22:@19747.4]
  assign dot_6_io_b_7 = $signed(io_wgt_data_bits_6_7); // @[TensorGemm.scala 165:22:@19751.4]
  assign dot_6_io_b_8 = $signed(io_wgt_data_bits_6_8); // @[TensorGemm.scala 165:22:@19755.4]
  assign dot_6_io_b_9 = $signed(io_wgt_data_bits_6_9); // @[TensorGemm.scala 165:22:@19759.4]
  assign dot_6_io_b_10 = $signed(io_wgt_data_bits_6_10); // @[TensorGemm.scala 165:22:@19763.4]
  assign dot_6_io_b_11 = $signed(io_wgt_data_bits_6_11); // @[TensorGemm.scala 165:22:@19767.4]
  assign dot_6_io_b_12 = $signed(io_wgt_data_bits_6_12); // @[TensorGemm.scala 165:22:@19771.4]
  assign dot_6_io_b_13 = $signed(io_wgt_data_bits_6_13); // @[TensorGemm.scala 165:22:@19775.4]
  assign dot_6_io_b_14 = $signed(io_wgt_data_bits_6_14); // @[TensorGemm.scala 165:22:@19779.4]
  assign dot_6_io_b_15 = $signed(io_wgt_data_bits_6_15); // @[TensorGemm.scala 165:22:@19783.4]
  assign dot_7_clock = clock; // @[:@19137.4]
  assign dot_7_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19802.4]
  assign dot_7_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19806.4]
  assign dot_7_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19810.4]
  assign dot_7_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19814.4]
  assign dot_7_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19818.4]
  assign dot_7_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19822.4]
  assign dot_7_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19826.4]
  assign dot_7_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19830.4]
  assign dot_7_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19834.4]
  assign dot_7_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19838.4]
  assign dot_7_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19842.4]
  assign dot_7_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19846.4]
  assign dot_7_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19850.4]
  assign dot_7_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19854.4]
  assign dot_7_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19858.4]
  assign dot_7_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19862.4]
  assign dot_7_io_b_0 = $signed(io_wgt_data_bits_7_0); // @[TensorGemm.scala 165:22:@19804.4]
  assign dot_7_io_b_1 = $signed(io_wgt_data_bits_7_1); // @[TensorGemm.scala 165:22:@19808.4]
  assign dot_7_io_b_2 = $signed(io_wgt_data_bits_7_2); // @[TensorGemm.scala 165:22:@19812.4]
  assign dot_7_io_b_3 = $signed(io_wgt_data_bits_7_3); // @[TensorGemm.scala 165:22:@19816.4]
  assign dot_7_io_b_4 = $signed(io_wgt_data_bits_7_4); // @[TensorGemm.scala 165:22:@19820.4]
  assign dot_7_io_b_5 = $signed(io_wgt_data_bits_7_5); // @[TensorGemm.scala 165:22:@19824.4]
  assign dot_7_io_b_6 = $signed(io_wgt_data_bits_7_6); // @[TensorGemm.scala 165:22:@19828.4]
  assign dot_7_io_b_7 = $signed(io_wgt_data_bits_7_7); // @[TensorGemm.scala 165:22:@19832.4]
  assign dot_7_io_b_8 = $signed(io_wgt_data_bits_7_8); // @[TensorGemm.scala 165:22:@19836.4]
  assign dot_7_io_b_9 = $signed(io_wgt_data_bits_7_9); // @[TensorGemm.scala 165:22:@19840.4]
  assign dot_7_io_b_10 = $signed(io_wgt_data_bits_7_10); // @[TensorGemm.scala 165:22:@19844.4]
  assign dot_7_io_b_11 = $signed(io_wgt_data_bits_7_11); // @[TensorGemm.scala 165:22:@19848.4]
  assign dot_7_io_b_12 = $signed(io_wgt_data_bits_7_12); // @[TensorGemm.scala 165:22:@19852.4]
  assign dot_7_io_b_13 = $signed(io_wgt_data_bits_7_13); // @[TensorGemm.scala 165:22:@19856.4]
  assign dot_7_io_b_14 = $signed(io_wgt_data_bits_7_14); // @[TensorGemm.scala 165:22:@19860.4]
  assign dot_7_io_b_15 = $signed(io_wgt_data_bits_7_15); // @[TensorGemm.scala 165:22:@19864.4]
  assign dot_8_clock = clock; // @[:@19140.4]
  assign dot_8_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19883.4]
  assign dot_8_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19887.4]
  assign dot_8_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19891.4]
  assign dot_8_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19895.4]
  assign dot_8_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19899.4]
  assign dot_8_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19903.4]
  assign dot_8_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19907.4]
  assign dot_8_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19911.4]
  assign dot_8_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19915.4]
  assign dot_8_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@19919.4]
  assign dot_8_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@19923.4]
  assign dot_8_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@19927.4]
  assign dot_8_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@19931.4]
  assign dot_8_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@19935.4]
  assign dot_8_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@19939.4]
  assign dot_8_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@19943.4]
  assign dot_8_io_b_0 = $signed(io_wgt_data_bits_8_0); // @[TensorGemm.scala 165:22:@19885.4]
  assign dot_8_io_b_1 = $signed(io_wgt_data_bits_8_1); // @[TensorGemm.scala 165:22:@19889.4]
  assign dot_8_io_b_2 = $signed(io_wgt_data_bits_8_2); // @[TensorGemm.scala 165:22:@19893.4]
  assign dot_8_io_b_3 = $signed(io_wgt_data_bits_8_3); // @[TensorGemm.scala 165:22:@19897.4]
  assign dot_8_io_b_4 = $signed(io_wgt_data_bits_8_4); // @[TensorGemm.scala 165:22:@19901.4]
  assign dot_8_io_b_5 = $signed(io_wgt_data_bits_8_5); // @[TensorGemm.scala 165:22:@19905.4]
  assign dot_8_io_b_6 = $signed(io_wgt_data_bits_8_6); // @[TensorGemm.scala 165:22:@19909.4]
  assign dot_8_io_b_7 = $signed(io_wgt_data_bits_8_7); // @[TensorGemm.scala 165:22:@19913.4]
  assign dot_8_io_b_8 = $signed(io_wgt_data_bits_8_8); // @[TensorGemm.scala 165:22:@19917.4]
  assign dot_8_io_b_9 = $signed(io_wgt_data_bits_8_9); // @[TensorGemm.scala 165:22:@19921.4]
  assign dot_8_io_b_10 = $signed(io_wgt_data_bits_8_10); // @[TensorGemm.scala 165:22:@19925.4]
  assign dot_8_io_b_11 = $signed(io_wgt_data_bits_8_11); // @[TensorGemm.scala 165:22:@19929.4]
  assign dot_8_io_b_12 = $signed(io_wgt_data_bits_8_12); // @[TensorGemm.scala 165:22:@19933.4]
  assign dot_8_io_b_13 = $signed(io_wgt_data_bits_8_13); // @[TensorGemm.scala 165:22:@19937.4]
  assign dot_8_io_b_14 = $signed(io_wgt_data_bits_8_14); // @[TensorGemm.scala 165:22:@19941.4]
  assign dot_8_io_b_15 = $signed(io_wgt_data_bits_8_15); // @[TensorGemm.scala 165:22:@19945.4]
  assign dot_9_clock = clock; // @[:@19143.4]
  assign dot_9_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@19964.4]
  assign dot_9_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@19968.4]
  assign dot_9_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@19972.4]
  assign dot_9_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@19976.4]
  assign dot_9_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@19980.4]
  assign dot_9_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@19984.4]
  assign dot_9_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@19988.4]
  assign dot_9_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@19992.4]
  assign dot_9_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@19996.4]
  assign dot_9_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@20000.4]
  assign dot_9_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@20004.4]
  assign dot_9_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@20008.4]
  assign dot_9_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@20012.4]
  assign dot_9_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@20016.4]
  assign dot_9_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@20020.4]
  assign dot_9_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@20024.4]
  assign dot_9_io_b_0 = $signed(io_wgt_data_bits_9_0); // @[TensorGemm.scala 165:22:@19966.4]
  assign dot_9_io_b_1 = $signed(io_wgt_data_bits_9_1); // @[TensorGemm.scala 165:22:@19970.4]
  assign dot_9_io_b_2 = $signed(io_wgt_data_bits_9_2); // @[TensorGemm.scala 165:22:@19974.4]
  assign dot_9_io_b_3 = $signed(io_wgt_data_bits_9_3); // @[TensorGemm.scala 165:22:@19978.4]
  assign dot_9_io_b_4 = $signed(io_wgt_data_bits_9_4); // @[TensorGemm.scala 165:22:@19982.4]
  assign dot_9_io_b_5 = $signed(io_wgt_data_bits_9_5); // @[TensorGemm.scala 165:22:@19986.4]
  assign dot_9_io_b_6 = $signed(io_wgt_data_bits_9_6); // @[TensorGemm.scala 165:22:@19990.4]
  assign dot_9_io_b_7 = $signed(io_wgt_data_bits_9_7); // @[TensorGemm.scala 165:22:@19994.4]
  assign dot_9_io_b_8 = $signed(io_wgt_data_bits_9_8); // @[TensorGemm.scala 165:22:@19998.4]
  assign dot_9_io_b_9 = $signed(io_wgt_data_bits_9_9); // @[TensorGemm.scala 165:22:@20002.4]
  assign dot_9_io_b_10 = $signed(io_wgt_data_bits_9_10); // @[TensorGemm.scala 165:22:@20006.4]
  assign dot_9_io_b_11 = $signed(io_wgt_data_bits_9_11); // @[TensorGemm.scala 165:22:@20010.4]
  assign dot_9_io_b_12 = $signed(io_wgt_data_bits_9_12); // @[TensorGemm.scala 165:22:@20014.4]
  assign dot_9_io_b_13 = $signed(io_wgt_data_bits_9_13); // @[TensorGemm.scala 165:22:@20018.4]
  assign dot_9_io_b_14 = $signed(io_wgt_data_bits_9_14); // @[TensorGemm.scala 165:22:@20022.4]
  assign dot_9_io_b_15 = $signed(io_wgt_data_bits_9_15); // @[TensorGemm.scala 165:22:@20026.4]
  assign dot_10_clock = clock; // @[:@19146.4]
  assign dot_10_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@20045.4]
  assign dot_10_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@20049.4]
  assign dot_10_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@20053.4]
  assign dot_10_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@20057.4]
  assign dot_10_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@20061.4]
  assign dot_10_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@20065.4]
  assign dot_10_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@20069.4]
  assign dot_10_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@20073.4]
  assign dot_10_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@20077.4]
  assign dot_10_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@20081.4]
  assign dot_10_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@20085.4]
  assign dot_10_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@20089.4]
  assign dot_10_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@20093.4]
  assign dot_10_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@20097.4]
  assign dot_10_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@20101.4]
  assign dot_10_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@20105.4]
  assign dot_10_io_b_0 = $signed(io_wgt_data_bits_10_0); // @[TensorGemm.scala 165:22:@20047.4]
  assign dot_10_io_b_1 = $signed(io_wgt_data_bits_10_1); // @[TensorGemm.scala 165:22:@20051.4]
  assign dot_10_io_b_2 = $signed(io_wgt_data_bits_10_2); // @[TensorGemm.scala 165:22:@20055.4]
  assign dot_10_io_b_3 = $signed(io_wgt_data_bits_10_3); // @[TensorGemm.scala 165:22:@20059.4]
  assign dot_10_io_b_4 = $signed(io_wgt_data_bits_10_4); // @[TensorGemm.scala 165:22:@20063.4]
  assign dot_10_io_b_5 = $signed(io_wgt_data_bits_10_5); // @[TensorGemm.scala 165:22:@20067.4]
  assign dot_10_io_b_6 = $signed(io_wgt_data_bits_10_6); // @[TensorGemm.scala 165:22:@20071.4]
  assign dot_10_io_b_7 = $signed(io_wgt_data_bits_10_7); // @[TensorGemm.scala 165:22:@20075.4]
  assign dot_10_io_b_8 = $signed(io_wgt_data_bits_10_8); // @[TensorGemm.scala 165:22:@20079.4]
  assign dot_10_io_b_9 = $signed(io_wgt_data_bits_10_9); // @[TensorGemm.scala 165:22:@20083.4]
  assign dot_10_io_b_10 = $signed(io_wgt_data_bits_10_10); // @[TensorGemm.scala 165:22:@20087.4]
  assign dot_10_io_b_11 = $signed(io_wgt_data_bits_10_11); // @[TensorGemm.scala 165:22:@20091.4]
  assign dot_10_io_b_12 = $signed(io_wgt_data_bits_10_12); // @[TensorGemm.scala 165:22:@20095.4]
  assign dot_10_io_b_13 = $signed(io_wgt_data_bits_10_13); // @[TensorGemm.scala 165:22:@20099.4]
  assign dot_10_io_b_14 = $signed(io_wgt_data_bits_10_14); // @[TensorGemm.scala 165:22:@20103.4]
  assign dot_10_io_b_15 = $signed(io_wgt_data_bits_10_15); // @[TensorGemm.scala 165:22:@20107.4]
  assign dot_11_clock = clock; // @[:@19149.4]
  assign dot_11_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@20126.4]
  assign dot_11_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@20130.4]
  assign dot_11_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@20134.4]
  assign dot_11_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@20138.4]
  assign dot_11_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@20142.4]
  assign dot_11_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@20146.4]
  assign dot_11_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@20150.4]
  assign dot_11_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@20154.4]
  assign dot_11_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@20158.4]
  assign dot_11_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@20162.4]
  assign dot_11_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@20166.4]
  assign dot_11_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@20170.4]
  assign dot_11_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@20174.4]
  assign dot_11_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@20178.4]
  assign dot_11_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@20182.4]
  assign dot_11_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@20186.4]
  assign dot_11_io_b_0 = $signed(io_wgt_data_bits_11_0); // @[TensorGemm.scala 165:22:@20128.4]
  assign dot_11_io_b_1 = $signed(io_wgt_data_bits_11_1); // @[TensorGemm.scala 165:22:@20132.4]
  assign dot_11_io_b_2 = $signed(io_wgt_data_bits_11_2); // @[TensorGemm.scala 165:22:@20136.4]
  assign dot_11_io_b_3 = $signed(io_wgt_data_bits_11_3); // @[TensorGemm.scala 165:22:@20140.4]
  assign dot_11_io_b_4 = $signed(io_wgt_data_bits_11_4); // @[TensorGemm.scala 165:22:@20144.4]
  assign dot_11_io_b_5 = $signed(io_wgt_data_bits_11_5); // @[TensorGemm.scala 165:22:@20148.4]
  assign dot_11_io_b_6 = $signed(io_wgt_data_bits_11_6); // @[TensorGemm.scala 165:22:@20152.4]
  assign dot_11_io_b_7 = $signed(io_wgt_data_bits_11_7); // @[TensorGemm.scala 165:22:@20156.4]
  assign dot_11_io_b_8 = $signed(io_wgt_data_bits_11_8); // @[TensorGemm.scala 165:22:@20160.4]
  assign dot_11_io_b_9 = $signed(io_wgt_data_bits_11_9); // @[TensorGemm.scala 165:22:@20164.4]
  assign dot_11_io_b_10 = $signed(io_wgt_data_bits_11_10); // @[TensorGemm.scala 165:22:@20168.4]
  assign dot_11_io_b_11 = $signed(io_wgt_data_bits_11_11); // @[TensorGemm.scala 165:22:@20172.4]
  assign dot_11_io_b_12 = $signed(io_wgt_data_bits_11_12); // @[TensorGemm.scala 165:22:@20176.4]
  assign dot_11_io_b_13 = $signed(io_wgt_data_bits_11_13); // @[TensorGemm.scala 165:22:@20180.4]
  assign dot_11_io_b_14 = $signed(io_wgt_data_bits_11_14); // @[TensorGemm.scala 165:22:@20184.4]
  assign dot_11_io_b_15 = $signed(io_wgt_data_bits_11_15); // @[TensorGemm.scala 165:22:@20188.4]
  assign dot_12_clock = clock; // @[:@19152.4]
  assign dot_12_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@20207.4]
  assign dot_12_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@20211.4]
  assign dot_12_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@20215.4]
  assign dot_12_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@20219.4]
  assign dot_12_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@20223.4]
  assign dot_12_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@20227.4]
  assign dot_12_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@20231.4]
  assign dot_12_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@20235.4]
  assign dot_12_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@20239.4]
  assign dot_12_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@20243.4]
  assign dot_12_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@20247.4]
  assign dot_12_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@20251.4]
  assign dot_12_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@20255.4]
  assign dot_12_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@20259.4]
  assign dot_12_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@20263.4]
  assign dot_12_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@20267.4]
  assign dot_12_io_b_0 = $signed(io_wgt_data_bits_12_0); // @[TensorGemm.scala 165:22:@20209.4]
  assign dot_12_io_b_1 = $signed(io_wgt_data_bits_12_1); // @[TensorGemm.scala 165:22:@20213.4]
  assign dot_12_io_b_2 = $signed(io_wgt_data_bits_12_2); // @[TensorGemm.scala 165:22:@20217.4]
  assign dot_12_io_b_3 = $signed(io_wgt_data_bits_12_3); // @[TensorGemm.scala 165:22:@20221.4]
  assign dot_12_io_b_4 = $signed(io_wgt_data_bits_12_4); // @[TensorGemm.scala 165:22:@20225.4]
  assign dot_12_io_b_5 = $signed(io_wgt_data_bits_12_5); // @[TensorGemm.scala 165:22:@20229.4]
  assign dot_12_io_b_6 = $signed(io_wgt_data_bits_12_6); // @[TensorGemm.scala 165:22:@20233.4]
  assign dot_12_io_b_7 = $signed(io_wgt_data_bits_12_7); // @[TensorGemm.scala 165:22:@20237.4]
  assign dot_12_io_b_8 = $signed(io_wgt_data_bits_12_8); // @[TensorGemm.scala 165:22:@20241.4]
  assign dot_12_io_b_9 = $signed(io_wgt_data_bits_12_9); // @[TensorGemm.scala 165:22:@20245.4]
  assign dot_12_io_b_10 = $signed(io_wgt_data_bits_12_10); // @[TensorGemm.scala 165:22:@20249.4]
  assign dot_12_io_b_11 = $signed(io_wgt_data_bits_12_11); // @[TensorGemm.scala 165:22:@20253.4]
  assign dot_12_io_b_12 = $signed(io_wgt_data_bits_12_12); // @[TensorGemm.scala 165:22:@20257.4]
  assign dot_12_io_b_13 = $signed(io_wgt_data_bits_12_13); // @[TensorGemm.scala 165:22:@20261.4]
  assign dot_12_io_b_14 = $signed(io_wgt_data_bits_12_14); // @[TensorGemm.scala 165:22:@20265.4]
  assign dot_12_io_b_15 = $signed(io_wgt_data_bits_12_15); // @[TensorGemm.scala 165:22:@20269.4]
  assign dot_13_clock = clock; // @[:@19155.4]
  assign dot_13_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@20288.4]
  assign dot_13_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@20292.4]
  assign dot_13_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@20296.4]
  assign dot_13_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@20300.4]
  assign dot_13_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@20304.4]
  assign dot_13_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@20308.4]
  assign dot_13_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@20312.4]
  assign dot_13_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@20316.4]
  assign dot_13_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@20320.4]
  assign dot_13_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@20324.4]
  assign dot_13_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@20328.4]
  assign dot_13_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@20332.4]
  assign dot_13_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@20336.4]
  assign dot_13_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@20340.4]
  assign dot_13_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@20344.4]
  assign dot_13_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@20348.4]
  assign dot_13_io_b_0 = $signed(io_wgt_data_bits_13_0); // @[TensorGemm.scala 165:22:@20290.4]
  assign dot_13_io_b_1 = $signed(io_wgt_data_bits_13_1); // @[TensorGemm.scala 165:22:@20294.4]
  assign dot_13_io_b_2 = $signed(io_wgt_data_bits_13_2); // @[TensorGemm.scala 165:22:@20298.4]
  assign dot_13_io_b_3 = $signed(io_wgt_data_bits_13_3); // @[TensorGemm.scala 165:22:@20302.4]
  assign dot_13_io_b_4 = $signed(io_wgt_data_bits_13_4); // @[TensorGemm.scala 165:22:@20306.4]
  assign dot_13_io_b_5 = $signed(io_wgt_data_bits_13_5); // @[TensorGemm.scala 165:22:@20310.4]
  assign dot_13_io_b_6 = $signed(io_wgt_data_bits_13_6); // @[TensorGemm.scala 165:22:@20314.4]
  assign dot_13_io_b_7 = $signed(io_wgt_data_bits_13_7); // @[TensorGemm.scala 165:22:@20318.4]
  assign dot_13_io_b_8 = $signed(io_wgt_data_bits_13_8); // @[TensorGemm.scala 165:22:@20322.4]
  assign dot_13_io_b_9 = $signed(io_wgt_data_bits_13_9); // @[TensorGemm.scala 165:22:@20326.4]
  assign dot_13_io_b_10 = $signed(io_wgt_data_bits_13_10); // @[TensorGemm.scala 165:22:@20330.4]
  assign dot_13_io_b_11 = $signed(io_wgt_data_bits_13_11); // @[TensorGemm.scala 165:22:@20334.4]
  assign dot_13_io_b_12 = $signed(io_wgt_data_bits_13_12); // @[TensorGemm.scala 165:22:@20338.4]
  assign dot_13_io_b_13 = $signed(io_wgt_data_bits_13_13); // @[TensorGemm.scala 165:22:@20342.4]
  assign dot_13_io_b_14 = $signed(io_wgt_data_bits_13_14); // @[TensorGemm.scala 165:22:@20346.4]
  assign dot_13_io_b_15 = $signed(io_wgt_data_bits_13_15); // @[TensorGemm.scala 165:22:@20350.4]
  assign dot_14_clock = clock; // @[:@19158.4]
  assign dot_14_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@20369.4]
  assign dot_14_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@20373.4]
  assign dot_14_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@20377.4]
  assign dot_14_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@20381.4]
  assign dot_14_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@20385.4]
  assign dot_14_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@20389.4]
  assign dot_14_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@20393.4]
  assign dot_14_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@20397.4]
  assign dot_14_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@20401.4]
  assign dot_14_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@20405.4]
  assign dot_14_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@20409.4]
  assign dot_14_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@20413.4]
  assign dot_14_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@20417.4]
  assign dot_14_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@20421.4]
  assign dot_14_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@20425.4]
  assign dot_14_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@20429.4]
  assign dot_14_io_b_0 = $signed(io_wgt_data_bits_14_0); // @[TensorGemm.scala 165:22:@20371.4]
  assign dot_14_io_b_1 = $signed(io_wgt_data_bits_14_1); // @[TensorGemm.scala 165:22:@20375.4]
  assign dot_14_io_b_2 = $signed(io_wgt_data_bits_14_2); // @[TensorGemm.scala 165:22:@20379.4]
  assign dot_14_io_b_3 = $signed(io_wgt_data_bits_14_3); // @[TensorGemm.scala 165:22:@20383.4]
  assign dot_14_io_b_4 = $signed(io_wgt_data_bits_14_4); // @[TensorGemm.scala 165:22:@20387.4]
  assign dot_14_io_b_5 = $signed(io_wgt_data_bits_14_5); // @[TensorGemm.scala 165:22:@20391.4]
  assign dot_14_io_b_6 = $signed(io_wgt_data_bits_14_6); // @[TensorGemm.scala 165:22:@20395.4]
  assign dot_14_io_b_7 = $signed(io_wgt_data_bits_14_7); // @[TensorGemm.scala 165:22:@20399.4]
  assign dot_14_io_b_8 = $signed(io_wgt_data_bits_14_8); // @[TensorGemm.scala 165:22:@20403.4]
  assign dot_14_io_b_9 = $signed(io_wgt_data_bits_14_9); // @[TensorGemm.scala 165:22:@20407.4]
  assign dot_14_io_b_10 = $signed(io_wgt_data_bits_14_10); // @[TensorGemm.scala 165:22:@20411.4]
  assign dot_14_io_b_11 = $signed(io_wgt_data_bits_14_11); // @[TensorGemm.scala 165:22:@20415.4]
  assign dot_14_io_b_12 = $signed(io_wgt_data_bits_14_12); // @[TensorGemm.scala 165:22:@20419.4]
  assign dot_14_io_b_13 = $signed(io_wgt_data_bits_14_13); // @[TensorGemm.scala 165:22:@20423.4]
  assign dot_14_io_b_14 = $signed(io_wgt_data_bits_14_14); // @[TensorGemm.scala 165:22:@20427.4]
  assign dot_14_io_b_15 = $signed(io_wgt_data_bits_14_15); // @[TensorGemm.scala 165:22:@20431.4]
  assign dot_15_clock = clock; // @[:@19161.4]
  assign dot_15_io_a_0 = $signed(io_inp_data_bits_0_0); // @[TensorGemm.scala 164:22:@20450.4]
  assign dot_15_io_a_1 = $signed(io_inp_data_bits_0_1); // @[TensorGemm.scala 164:22:@20454.4]
  assign dot_15_io_a_2 = $signed(io_inp_data_bits_0_2); // @[TensorGemm.scala 164:22:@20458.4]
  assign dot_15_io_a_3 = $signed(io_inp_data_bits_0_3); // @[TensorGemm.scala 164:22:@20462.4]
  assign dot_15_io_a_4 = $signed(io_inp_data_bits_0_4); // @[TensorGemm.scala 164:22:@20466.4]
  assign dot_15_io_a_5 = $signed(io_inp_data_bits_0_5); // @[TensorGemm.scala 164:22:@20470.4]
  assign dot_15_io_a_6 = $signed(io_inp_data_bits_0_6); // @[TensorGemm.scala 164:22:@20474.4]
  assign dot_15_io_a_7 = $signed(io_inp_data_bits_0_7); // @[TensorGemm.scala 164:22:@20478.4]
  assign dot_15_io_a_8 = $signed(io_inp_data_bits_0_8); // @[TensorGemm.scala 164:22:@20482.4]
  assign dot_15_io_a_9 = $signed(io_inp_data_bits_0_9); // @[TensorGemm.scala 164:22:@20486.4]
  assign dot_15_io_a_10 = $signed(io_inp_data_bits_0_10); // @[TensorGemm.scala 164:22:@20490.4]
  assign dot_15_io_a_11 = $signed(io_inp_data_bits_0_11); // @[TensorGemm.scala 164:22:@20494.4]
  assign dot_15_io_a_12 = $signed(io_inp_data_bits_0_12); // @[TensorGemm.scala 164:22:@20498.4]
  assign dot_15_io_a_13 = $signed(io_inp_data_bits_0_13); // @[TensorGemm.scala 164:22:@20502.4]
  assign dot_15_io_a_14 = $signed(io_inp_data_bits_0_14); // @[TensorGemm.scala 164:22:@20506.4]
  assign dot_15_io_a_15 = $signed(io_inp_data_bits_0_15); // @[TensorGemm.scala 164:22:@20510.4]
  assign dot_15_io_b_0 = $signed(io_wgt_data_bits_15_0); // @[TensorGemm.scala 165:22:@20452.4]
  assign dot_15_io_b_1 = $signed(io_wgt_data_bits_15_1); // @[TensorGemm.scala 165:22:@20456.4]
  assign dot_15_io_b_2 = $signed(io_wgt_data_bits_15_2); // @[TensorGemm.scala 165:22:@20460.4]
  assign dot_15_io_b_3 = $signed(io_wgt_data_bits_15_3); // @[TensorGemm.scala 165:22:@20464.4]
  assign dot_15_io_b_4 = $signed(io_wgt_data_bits_15_4); // @[TensorGemm.scala 165:22:@20468.4]
  assign dot_15_io_b_5 = $signed(io_wgt_data_bits_15_5); // @[TensorGemm.scala 165:22:@20472.4]
  assign dot_15_io_b_6 = $signed(io_wgt_data_bits_15_6); // @[TensorGemm.scala 165:22:@20476.4]
  assign dot_15_io_b_7 = $signed(io_wgt_data_bits_15_7); // @[TensorGemm.scala 165:22:@20480.4]
  assign dot_15_io_b_8 = $signed(io_wgt_data_bits_15_8); // @[TensorGemm.scala 165:22:@20484.4]
  assign dot_15_io_b_9 = $signed(io_wgt_data_bits_15_9); // @[TensorGemm.scala 165:22:@20488.4]
  assign dot_15_io_b_10 = $signed(io_wgt_data_bits_15_10); // @[TensorGemm.scala 165:22:@20492.4]
  assign dot_15_io_b_11 = $signed(io_wgt_data_bits_15_11); // @[TensorGemm.scala 165:22:@20496.4]
  assign dot_15_io_b_12 = $signed(io_wgt_data_bits_15_12); // @[TensorGemm.scala 165:22:@20500.4]
  assign dot_15_io_b_13 = $signed(io_wgt_data_bits_15_13); // @[TensorGemm.scala 165:22:@20504.4]
  assign dot_15_io_b_14 = $signed(io_wgt_data_bits_15_14); // @[TensorGemm.scala 165:22:@20508.4]
  assign dot_15_io_b_15 = $signed(io_wgt_data_bits_15_15); // @[TensorGemm.scala 165:22:@20512.4]
  assign acc_0_clock = clock; // @[:@19164.4]
  assign acc_0_reset = reset; // @[:@19165.4]
  assign acc_0_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19232.4]
  assign acc_0_io_enq_bits = io_acc_i_data_bits_0_0; // @[TensorGemm.scala 162:24:@19233.4]
  assign acc_1_clock = clock; // @[:@19167.4]
  assign acc_1_reset = reset; // @[:@19168.4]
  assign acc_1_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19313.4]
  assign acc_1_io_enq_bits = io_acc_i_data_bits_0_1; // @[TensorGemm.scala 162:24:@19314.4]
  assign acc_2_clock = clock; // @[:@19170.4]
  assign acc_2_reset = reset; // @[:@19171.4]
  assign acc_2_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19394.4]
  assign acc_2_io_enq_bits = io_acc_i_data_bits_0_2; // @[TensorGemm.scala 162:24:@19395.4]
  assign acc_3_clock = clock; // @[:@19173.4]
  assign acc_3_reset = reset; // @[:@19174.4]
  assign acc_3_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19475.4]
  assign acc_3_io_enq_bits = io_acc_i_data_bits_0_3; // @[TensorGemm.scala 162:24:@19476.4]
  assign acc_4_clock = clock; // @[:@19176.4]
  assign acc_4_reset = reset; // @[:@19177.4]
  assign acc_4_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19556.4]
  assign acc_4_io_enq_bits = io_acc_i_data_bits_0_4; // @[TensorGemm.scala 162:24:@19557.4]
  assign acc_5_clock = clock; // @[:@19179.4]
  assign acc_5_reset = reset; // @[:@19180.4]
  assign acc_5_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19637.4]
  assign acc_5_io_enq_bits = io_acc_i_data_bits_0_5; // @[TensorGemm.scala 162:24:@19638.4]
  assign acc_6_clock = clock; // @[:@19182.4]
  assign acc_6_reset = reset; // @[:@19183.4]
  assign acc_6_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19718.4]
  assign acc_6_io_enq_bits = io_acc_i_data_bits_0_6; // @[TensorGemm.scala 162:24:@19719.4]
  assign acc_7_clock = clock; // @[:@19185.4]
  assign acc_7_reset = reset; // @[:@19186.4]
  assign acc_7_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19799.4]
  assign acc_7_io_enq_bits = io_acc_i_data_bits_0_7; // @[TensorGemm.scala 162:24:@19800.4]
  assign acc_8_clock = clock; // @[:@19188.4]
  assign acc_8_reset = reset; // @[:@19189.4]
  assign acc_8_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19880.4]
  assign acc_8_io_enq_bits = io_acc_i_data_bits_0_8; // @[TensorGemm.scala 162:24:@19881.4]
  assign acc_9_clock = clock; // @[:@19191.4]
  assign acc_9_reset = reset; // @[:@19192.4]
  assign acc_9_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@19961.4]
  assign acc_9_io_enq_bits = io_acc_i_data_bits_0_9; // @[TensorGemm.scala 162:24:@19962.4]
  assign acc_10_clock = clock; // @[:@19194.4]
  assign acc_10_reset = reset; // @[:@19195.4]
  assign acc_10_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@20042.4]
  assign acc_10_io_enq_bits = io_acc_i_data_bits_0_10; // @[TensorGemm.scala 162:24:@20043.4]
  assign acc_11_clock = clock; // @[:@19197.4]
  assign acc_11_reset = reset; // @[:@19198.4]
  assign acc_11_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@20123.4]
  assign acc_11_io_enq_bits = io_acc_i_data_bits_0_11; // @[TensorGemm.scala 162:24:@20124.4]
  assign acc_12_clock = clock; // @[:@19200.4]
  assign acc_12_reset = reset; // @[:@19201.4]
  assign acc_12_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@20204.4]
  assign acc_12_io_enq_bits = io_acc_i_data_bits_0_12; // @[TensorGemm.scala 162:24:@20205.4]
  assign acc_13_clock = clock; // @[:@19203.4]
  assign acc_13_reset = reset; // @[:@19204.4]
  assign acc_13_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@20285.4]
  assign acc_13_io_enq_bits = io_acc_i_data_bits_0_13; // @[TensorGemm.scala 162:24:@20286.4]
  assign acc_14_clock = clock; // @[:@19206.4]
  assign acc_14_reset = reset; // @[:@19207.4]
  assign acc_14_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@20366.4]
  assign acc_14_io_enq_bits = io_acc_i_data_bits_0_14; // @[TensorGemm.scala 162:24:@20367.4]
  assign acc_15_clock = clock; // @[:@19209.4]
  assign acc_15_reset = reset; // @[:@19210.4]
  assign acc_15_io_enq_valid = _T_6017 & _T_6018; // @[TensorGemm.scala 161:25:@20447.4]
  assign acc_15_io_enq_bits = io_acc_i_data_bits_0_15; // @[TensorGemm.scala 162:24:@20448.4]
endmodule
module Pipe_16( // @[:@20562.2]
  input         clock, // @[:@20563.4]
  input         reset, // @[:@20564.4]
  input         io_enq_valid, // @[:@20565.4]
  input  [13:0] io_enq_bits, // @[:@20565.4]
  output        io_deq_valid, // @[:@20565.4]
  output [13:0] io_deq_bits // @[:@20565.4]
);
  reg  _T_19; // @[Valid.scala 48:22:@20567.4]
  reg [31:0] _RAND_0;
  reg [13:0] _T_21; // @[Reg.scala 11:16:@20569.4]
  reg [31:0] _RAND_1;
  reg  _T_24; // @[Valid.scala 48:22:@20573.4]
  reg [31:0] _RAND_2;
  reg [13:0] _T_26; // @[Reg.scala 11:16:@20575.4]
  reg [31:0] _RAND_3;
  assign io_deq_valid = _T_24; // @[Valid.scala 70:10:@20583.4]
  assign io_deq_bits = _T_26; // @[Valid.scala 70:10:@20582.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_21 = _RAND_1[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_24 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_26 = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      _T_19 <= io_enq_valid;
    end
    if (io_enq_valid) begin
      _T_21 <= io_enq_bits;
    end
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_19;
    end
    if (_T_19) begin
      _T_26 <= _T_21;
    end
  end
endmodule
module TensorGemm( // @[:@20585.2]
  input          clock, // @[:@20586.4]
  input          reset, // @[:@20587.4]
  input          io_start, // @[:@20588.4]
  output         io_done, // @[:@20588.4]
  input  [127:0] io_inst, // @[:@20588.4]
  output         io_uop_idx_valid, // @[:@20588.4]
  output [10:0]  io_uop_idx_bits, // @[:@20588.4]
  input          io_uop_data_valid, // @[:@20588.4]
  input  [9:0]   io_uop_data_bits_u2, // @[:@20588.4]
  input  [10:0]  io_uop_data_bits_u1, // @[:@20588.4]
  input  [10:0]  io_uop_data_bits_u0, // @[:@20588.4]
  output         io_inp_rd_idx_valid, // @[:@20588.4]
  output [10:0]  io_inp_rd_idx_bits, // @[:@20588.4]
  input          io_inp_rd_data_valid, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_0, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_1, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_2, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_3, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_4, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_5, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_6, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_7, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_8, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_9, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_10, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_11, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_12, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_13, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_14, // @[:@20588.4]
  input  [7:0]   io_inp_rd_data_bits_0_15, // @[:@20588.4]
  output         io_wgt_rd_idx_valid, // @[:@20588.4]
  output [9:0]   io_wgt_rd_idx_bits, // @[:@20588.4]
  input          io_wgt_rd_data_valid, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_0_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_1_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_2_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_3_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_4_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_5_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_6_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_7_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_8_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_9_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_10_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_11_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_12_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_13_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_14_15, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_0, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_1, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_2, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_3, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_4, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_5, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_6, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_7, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_8, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_9, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_10, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_11, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_12, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_13, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_14, // @[:@20588.4]
  input  [7:0]   io_wgt_rd_data_bits_15_15, // @[:@20588.4]
  output         io_acc_rd_idx_valid, // @[:@20588.4]
  output [10:0]  io_acc_rd_idx_bits, // @[:@20588.4]
  input          io_acc_rd_data_valid, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_0, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_1, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_2, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_3, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_4, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_5, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_6, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_7, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_8, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_9, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_10, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_11, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_12, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_13, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_14, // @[:@20588.4]
  input  [31:0]  io_acc_rd_data_bits_0_15, // @[:@20588.4]
  output         io_acc_wr_valid, // @[:@20588.4]
  output [10:0]  io_acc_wr_bits_idx, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_0, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_1, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_2, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_3, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_4, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_5, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_6, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_7, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_8, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_9, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_10, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_11, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_12, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_13, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_14, // @[:@20588.4]
  output [31:0]  io_acc_wr_bits_data_0_15, // @[:@20588.4]
  output         io_out_wr_valid, // @[:@20588.4]
  output [10:0]  io_out_wr_bits_idx, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_0, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_1, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_2, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_3, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_4, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_5, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_6, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_7, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_8, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_9, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_10, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_11, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_12, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_13, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_14, // @[:@20588.4]
  output [7:0]   io_out_wr_bits_data_0_15 // @[:@20588.4]
);
  wire  mvc_clock; // @[TensorGemm.scala 199:19:@20591.4]
  wire  mvc_reset; // @[TensorGemm.scala 199:19:@20591.4]
  wire  mvc_io_reset; // @[TensorGemm.scala 199:19:@20591.4]
  wire  mvc_io_inp_data_valid; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_inp_data_bits_0_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire  mvc_io_wgt_data_valid; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_0_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_1_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_2_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_3_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_4_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_5_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_6_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_7_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_8_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_9_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_10_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_11_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_12_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_13_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_14_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_wgt_data_bits_15_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire  mvc_io_acc_i_data_valid; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_i_data_bits_0_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire  mvc_io_acc_o_data_valid; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [31:0] mvc_io_acc_o_data_bits_0_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire  mvc_io_out_data_valid; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_0; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_1; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_2; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_3; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_4; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_5; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_6; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_7; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_8; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_9; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_10; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_11; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_12; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_13; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_14; // @[TensorGemm.scala 199:19:@20591.4]
  wire [7:0] mvc_io_out_data_bits_0_15; // @[TensorGemm.scala 199:19:@20591.4]
  wire  wrpipe_clock; // @[TensorGemm.scala 218:22:@20644.4]
  wire  wrpipe_reset; // @[TensorGemm.scala 218:22:@20644.4]
  wire  wrpipe_io_enq_valid; // @[TensorGemm.scala 218:22:@20644.4]
  wire [13:0] wrpipe_io_enq_bits; // @[TensorGemm.scala 218:22:@20644.4]
  wire  wrpipe_io_deq_valid; // @[TensorGemm.scala 218:22:@20644.4]
  wire [13:0] wrpipe_io_deq_bits; // @[TensorGemm.scala 218:22:@20644.4]
  reg [2:0] state; // @[TensorGemm.scala 198:22:@20590.4]
  reg [31:0] _RAND_0;
  wire  dec_reset; // @[TensorGemm.scala 200:29:@20607.4]
  wire [12:0] dec_uop_begin; // @[TensorGemm.scala 200:29:@20609.4]
  wire [13:0] dec_uop_end; // @[TensorGemm.scala 200:29:@20611.4]
  wire [13:0] dec_lp_0; // @[TensorGemm.scala 200:29:@20613.4]
  wire [13:0] dec_lp_1; // @[TensorGemm.scala 200:29:@20615.4]
  wire [10:0] dec_acc_0; // @[TensorGemm.scala 200:29:@20619.4]
  wire [10:0] dec_acc_1; // @[TensorGemm.scala 200:29:@20621.4]
  wire [10:0] dec_inp_0; // @[TensorGemm.scala 200:29:@20623.4]
  wire [10:0] dec_inp_1; // @[TensorGemm.scala 200:29:@20625.4]
  wire [9:0] dec_wgt_0; // @[TensorGemm.scala 200:29:@20627.4]
  wire [9:0] dec_wgt_1; // @[TensorGemm.scala 200:29:@20629.4]
  reg [13:0] uop_idx; // @[TensorGemm.scala 201:20:@20631.4]
  reg [31:0] _RAND_1;
  reg [13:0] uop_acc; // @[TensorGemm.scala 203:20:@20632.4]
  reg [31:0] _RAND_2;
  reg [13:0] uop_inp; // @[TensorGemm.scala 204:20:@20633.4]
  reg [31:0] _RAND_3;
  reg [13:0] uop_wgt; // @[TensorGemm.scala 205:20:@20634.4]
  reg [31:0] _RAND_4;
  reg [13:0] cnt_o; // @[TensorGemm.scala 206:18:@20635.4]
  reg [31:0] _RAND_5;
  reg [13:0] acc_o; // @[TensorGemm.scala 207:18:@20636.4]
  reg [31:0] _RAND_6;
  reg [13:0] inp_o; // @[TensorGemm.scala 208:18:@20637.4]
  reg [31:0] _RAND_7;
  reg [13:0] wgt_o; // @[TensorGemm.scala 209:18:@20638.4]
  reg [31:0] _RAND_8;
  reg [13:0] cnt_i; // @[TensorGemm.scala 210:18:@20639.4]
  reg [31:0] _RAND_9;
  reg [13:0] acc_i; // @[TensorGemm.scala 211:18:@20640.4]
  reg [31:0] _RAND_10;
  reg [13:0] inp_i; // @[TensorGemm.scala 212:18:@20641.4]
  reg [31:0] _RAND_11;
  reg [13:0] wgt_i; // @[TensorGemm.scala 213:18:@20642.4]
  reg [31:0] _RAND_12;
  reg [4:0] inflight; // @[TensorGemm.scala 215:21:@20643.4]
  reg [31:0] _RAND_13;
  wire  _T_7688; // @[TensorGemm.scala 219:23:@20647.4]
  wire  _T_7689; // @[TensorGemm.scala 220:13:@20648.4]
  wire [14:0] _T_7691; // @[TensorGemm.scala 221:26:@20649.4]
  wire [14:0] _T_7692; // @[TensorGemm.scala 221:26:@20650.4]
  wire [13:0] _T_7693; // @[TensorGemm.scala 221:26:@20651.4]
  wire  _T_7694; // @[TensorGemm.scala 221:13:@20652.4]
  wire  _T_7695; // @[TensorGemm.scala 220:22:@20653.4]
  wire [14:0] _T_7697; // @[TensorGemm.scala 222:26:@20654.4]
  wire [14:0] _T_7698; // @[TensorGemm.scala 222:26:@20655.4]
  wire [13:0] _T_7699; // @[TensorGemm.scala 222:26:@20656.4]
  wire  _T_7700; // @[TensorGemm.scala 222:13:@20657.4]
  wire  _T_7701; // @[TensorGemm.scala 221:32:@20658.4]
  wire [14:0] _T_7703; // @[TensorGemm.scala 223:27:@20659.4]
  wire [14:0] _T_7704; // @[TensorGemm.scala 223:27:@20660.4]
  wire [13:0] _T_7705; // @[TensorGemm.scala 223:27:@20661.4]
  wire  _T_7706; // @[TensorGemm.scala 223:15:@20662.4]
  wire  _T_7707; // @[TensorGemm.scala 222:32:@20663.4]
  wire  _T_7710; // @[TensorGemm.scala 223:33:@20665.4]
  wire  _T_7711; // @[TensorGemm.scala 225:13:@20666.4]
  wire  _T_7712; // @[TensorGemm.scala 224:25:@20667.4]
  wire  _T_7713; // @[Conditional.scala 37:30:@20669.4]
  wire [2:0] _GEN_0; // @[TensorGemm.scala 229:22:@20671.6]
  wire  _T_7714; // @[Conditional.scala 37:30:@20676.6]
  wire  _T_7715; // @[Conditional.scala 37:30:@20681.8]
  wire  _T_7716; // @[Conditional.scala 37:30:@20686.10]
  wire  _T_7717; // @[Conditional.scala 37:30:@20691.12]
  wire  _T_7728; // @[TensorGemm.scala 244:36:@20701.14]
  wire  _T_7734; // @[TensorGemm.scala 245:38:@20706.14]
  wire  _T_7736; // @[TensorGemm.scala 247:23:@20708.16]
  wire [2:0] _GEN_1; // @[TensorGemm.scala 247:32:@20709.16]
  wire [2:0] _GEN_2; // @[TensorGemm.scala 246:40:@20707.14]
  wire  _T_7737; // @[Conditional.scala 37:30:@20721.14]
  wire [2:0] _GEN_3; // @[TensorGemm.scala 257:30:@20724.16]
  wire [2:0] _GEN_4; // @[Conditional.scala 39:67:@20722.14]
  wire [2:0] _GEN_5; // @[Conditional.scala 39:67:@20692.12]
  wire [2:0] _GEN_6; // @[Conditional.scala 39:67:@20687.10]
  wire [2:0] _GEN_7; // @[Conditional.scala 39:67:@20682.8]
  wire [2:0] _GEN_8; // @[Conditional.scala 39:67:@20677.6]
  wire [2:0] _GEN_9; // @[Conditional.scala 40:58:@20670.4]
  wire  _T_7740; // @[TensorGemm.scala 263:14:@20728.4]
  wire  _T_7743; // @[TensorGemm.scala 265:14:@20733.6]
  wire  _T_7744; // @[TensorGemm.scala 266:17:@20735.8]
  wire  _T_7745; // @[TensorGemm.scala 266:34:@20736.8]
  wire [5:0] _T_7748; // @[TensorGemm.scala 269:28:@20743.12]
  wire [4:0] _T_7749; // @[TensorGemm.scala 269:28:@20744.12]
  wire [5:0] _T_7751; // @[TensorGemm.scala 271:28:@20749.14]
  wire [5:0] _T_7752; // @[TensorGemm.scala 271:28:@20750.14]
  wire [4:0] _T_7753; // @[TensorGemm.scala 271:28:@20751.14]
  wire [4:0] _GEN_10; // @[TensorGemm.scala 270:41:@20748.12]
  wire [4:0] _GEN_11; // @[TensorGemm.scala 268:39:@20742.10]
  wire [4:0] _GEN_12; // @[TensorGemm.scala 266:62:@20737.8]
  wire [4:0] _GEN_13; // @[TensorGemm.scala 265:26:@20734.6]
  wire  _T_7761; // @[TensorGemm.scala 277:23:@20761.4]
  wire  _T_7762; // @[TensorGemm.scala 276:21:@20762.4]
  wire [13:0] _GEN_40; // @[TensorGemm.scala 280:46:@20768.6]
  wire  _T_7764; // @[TensorGemm.scala 280:46:@20768.6]
  wire  _T_7765; // @[TensorGemm.scala 280:29:@20769.6]
  wire [14:0] _T_7767; // @[TensorGemm.scala 281:24:@20771.8]
  wire [13:0] _T_7768; // @[TensorGemm.scala 281:24:@20772.8]
  wire [13:0] _GEN_15; // @[TensorGemm.scala 280:59:@20770.6]
  wire  _T_7786; // @[TensorGemm.scala 291:33:@20793.6]
  wire [14:0] _T_7788; // @[TensorGemm.scala 293:20:@20795.8]
  wire [13:0] _T_7789; // @[TensorGemm.scala 293:20:@20796.8]
  wire [13:0] _GEN_41; // @[TensorGemm.scala 294:20:@20798.8]
  wire [14:0] _T_7790; // @[TensorGemm.scala 294:20:@20798.8]
  wire [13:0] _T_7791; // @[TensorGemm.scala 294:20:@20799.8]
  wire [13:0] _GEN_42; // @[TensorGemm.scala 295:20:@20801.8]
  wire [14:0] _T_7792; // @[TensorGemm.scala 295:20:@20801.8]
  wire [13:0] _T_7793; // @[TensorGemm.scala 295:20:@20802.8]
  wire [13:0] _GEN_43; // @[TensorGemm.scala 296:20:@20804.8]
  wire [14:0] _T_7794; // @[TensorGemm.scala 296:20:@20804.8]
  wire [13:0] _T_7795; // @[TensorGemm.scala 296:20:@20805.8]
  wire [13:0] _GEN_17; // @[TensorGemm.scala 292:33:@20794.6]
  wire [13:0] _GEN_18; // @[TensorGemm.scala 292:33:@20794.6]
  wire [13:0] _GEN_19; // @[TensorGemm.scala 292:33:@20794.6]
  wire [13:0] _GEN_20; // @[TensorGemm.scala 292:33:@20794.6]
  wire  _T_7801; // @[TensorGemm.scala 304:20:@20816.6]
  wire  _T_7802; // @[TensorGemm.scala 304:42:@20817.6]
  wire  _T_7803; // @[TensorGemm.scala 304:33:@20818.6]
  wire [14:0] _T_7813; // @[TensorGemm.scala 310:20:@20833.10]
  wire [13:0] _T_7814; // @[TensorGemm.scala 310:20:@20834.10]
  wire [13:0] _GEN_44; // @[TensorGemm.scala 311:20:@20836.10]
  wire [14:0] _T_7815; // @[TensorGemm.scala 311:20:@20836.10]
  wire [13:0] _T_7816; // @[TensorGemm.scala 311:20:@20837.10]
  wire [13:0] _GEN_45; // @[TensorGemm.scala 312:20:@20839.10]
  wire [14:0] _T_7817; // @[TensorGemm.scala 312:20:@20839.10]
  wire [13:0] _T_7818; // @[TensorGemm.scala 312:20:@20840.10]
  wire [13:0] _GEN_46; // @[TensorGemm.scala 313:20:@20842.10]
  wire [14:0] _T_7819; // @[TensorGemm.scala 313:20:@20842.10]
  wire [13:0] _T_7820; // @[TensorGemm.scala 313:20:@20843.10]
  wire [13:0] _GEN_25; // @[TensorGemm.scala 309:59:@20832.8]
  wire [13:0] _GEN_26; // @[TensorGemm.scala 309:59:@20832.8]
  wire [13:0] _GEN_27; // @[TensorGemm.scala 309:59:@20832.8]
  wire [13:0] _GEN_28; // @[TensorGemm.scala 309:59:@20832.8]
  wire [13:0] _GEN_29; // @[TensorGemm.scala 304:56:@20819.6]
  wire [13:0] _GEN_30; // @[TensorGemm.scala 304:56:@20819.6]
  wire [13:0] _GEN_31; // @[TensorGemm.scala 304:56:@20819.6]
  wire [13:0] _GEN_32; // @[TensorGemm.scala 304:56:@20819.6]
  wire  _T_7821; // @[TensorGemm.scala 316:14:@20846.4]
  wire  _T_7822; // @[TensorGemm.scala 316:30:@20847.4]
  wire [13:0] _GEN_47; // @[TensorGemm.scala 317:36:@20849.6]
  wire [14:0] _T_7823; // @[TensorGemm.scala 317:36:@20849.6]
  wire [13:0] _T_7824; // @[TensorGemm.scala 317:36:@20850.6]
  wire [13:0] _GEN_48; // @[TensorGemm.scala 318:36:@20852.6]
  wire [14:0] _T_7825; // @[TensorGemm.scala 318:36:@20852.6]
  wire [13:0] _T_7826; // @[TensorGemm.scala 318:36:@20853.6]
  wire [13:0] _GEN_49; // @[TensorGemm.scala 319:36:@20855.6]
  wire [14:0] _T_7827; // @[TensorGemm.scala 319:36:@20855.6]
  wire [13:0] _T_7828; // @[TensorGemm.scala 319:36:@20856.6]
  wire  _T_7830; // @[TensorGemm.scala 322:43:@20860.4]
  wire  _T_8115; // @[TensorGemm.scala 351:8:@21446.4]
  wire [13:0] _T_8117; // @[TensorGemm.scala 352:28:@21449.4]
  MatrixVectorMultiplication mvc ( // @[TensorGemm.scala 199:19:@20591.4]
    .clock(mvc_clock),
    .reset(mvc_reset),
    .io_reset(mvc_io_reset),
    .io_inp_data_valid(mvc_io_inp_data_valid),
    .io_inp_data_bits_0_0(mvc_io_inp_data_bits_0_0),
    .io_inp_data_bits_0_1(mvc_io_inp_data_bits_0_1),
    .io_inp_data_bits_0_2(mvc_io_inp_data_bits_0_2),
    .io_inp_data_bits_0_3(mvc_io_inp_data_bits_0_3),
    .io_inp_data_bits_0_4(mvc_io_inp_data_bits_0_4),
    .io_inp_data_bits_0_5(mvc_io_inp_data_bits_0_5),
    .io_inp_data_bits_0_6(mvc_io_inp_data_bits_0_6),
    .io_inp_data_bits_0_7(mvc_io_inp_data_bits_0_7),
    .io_inp_data_bits_0_8(mvc_io_inp_data_bits_0_8),
    .io_inp_data_bits_0_9(mvc_io_inp_data_bits_0_9),
    .io_inp_data_bits_0_10(mvc_io_inp_data_bits_0_10),
    .io_inp_data_bits_0_11(mvc_io_inp_data_bits_0_11),
    .io_inp_data_bits_0_12(mvc_io_inp_data_bits_0_12),
    .io_inp_data_bits_0_13(mvc_io_inp_data_bits_0_13),
    .io_inp_data_bits_0_14(mvc_io_inp_data_bits_0_14),
    .io_inp_data_bits_0_15(mvc_io_inp_data_bits_0_15),
    .io_wgt_data_valid(mvc_io_wgt_data_valid),
    .io_wgt_data_bits_0_0(mvc_io_wgt_data_bits_0_0),
    .io_wgt_data_bits_0_1(mvc_io_wgt_data_bits_0_1),
    .io_wgt_data_bits_0_2(mvc_io_wgt_data_bits_0_2),
    .io_wgt_data_bits_0_3(mvc_io_wgt_data_bits_0_3),
    .io_wgt_data_bits_0_4(mvc_io_wgt_data_bits_0_4),
    .io_wgt_data_bits_0_5(mvc_io_wgt_data_bits_0_5),
    .io_wgt_data_bits_0_6(mvc_io_wgt_data_bits_0_6),
    .io_wgt_data_bits_0_7(mvc_io_wgt_data_bits_0_7),
    .io_wgt_data_bits_0_8(mvc_io_wgt_data_bits_0_8),
    .io_wgt_data_bits_0_9(mvc_io_wgt_data_bits_0_9),
    .io_wgt_data_bits_0_10(mvc_io_wgt_data_bits_0_10),
    .io_wgt_data_bits_0_11(mvc_io_wgt_data_bits_0_11),
    .io_wgt_data_bits_0_12(mvc_io_wgt_data_bits_0_12),
    .io_wgt_data_bits_0_13(mvc_io_wgt_data_bits_0_13),
    .io_wgt_data_bits_0_14(mvc_io_wgt_data_bits_0_14),
    .io_wgt_data_bits_0_15(mvc_io_wgt_data_bits_0_15),
    .io_wgt_data_bits_1_0(mvc_io_wgt_data_bits_1_0),
    .io_wgt_data_bits_1_1(mvc_io_wgt_data_bits_1_1),
    .io_wgt_data_bits_1_2(mvc_io_wgt_data_bits_1_2),
    .io_wgt_data_bits_1_3(mvc_io_wgt_data_bits_1_3),
    .io_wgt_data_bits_1_4(mvc_io_wgt_data_bits_1_4),
    .io_wgt_data_bits_1_5(mvc_io_wgt_data_bits_1_5),
    .io_wgt_data_bits_1_6(mvc_io_wgt_data_bits_1_6),
    .io_wgt_data_bits_1_7(mvc_io_wgt_data_bits_1_7),
    .io_wgt_data_bits_1_8(mvc_io_wgt_data_bits_1_8),
    .io_wgt_data_bits_1_9(mvc_io_wgt_data_bits_1_9),
    .io_wgt_data_bits_1_10(mvc_io_wgt_data_bits_1_10),
    .io_wgt_data_bits_1_11(mvc_io_wgt_data_bits_1_11),
    .io_wgt_data_bits_1_12(mvc_io_wgt_data_bits_1_12),
    .io_wgt_data_bits_1_13(mvc_io_wgt_data_bits_1_13),
    .io_wgt_data_bits_1_14(mvc_io_wgt_data_bits_1_14),
    .io_wgt_data_bits_1_15(mvc_io_wgt_data_bits_1_15),
    .io_wgt_data_bits_2_0(mvc_io_wgt_data_bits_2_0),
    .io_wgt_data_bits_2_1(mvc_io_wgt_data_bits_2_1),
    .io_wgt_data_bits_2_2(mvc_io_wgt_data_bits_2_2),
    .io_wgt_data_bits_2_3(mvc_io_wgt_data_bits_2_3),
    .io_wgt_data_bits_2_4(mvc_io_wgt_data_bits_2_4),
    .io_wgt_data_bits_2_5(mvc_io_wgt_data_bits_2_5),
    .io_wgt_data_bits_2_6(mvc_io_wgt_data_bits_2_6),
    .io_wgt_data_bits_2_7(mvc_io_wgt_data_bits_2_7),
    .io_wgt_data_bits_2_8(mvc_io_wgt_data_bits_2_8),
    .io_wgt_data_bits_2_9(mvc_io_wgt_data_bits_2_9),
    .io_wgt_data_bits_2_10(mvc_io_wgt_data_bits_2_10),
    .io_wgt_data_bits_2_11(mvc_io_wgt_data_bits_2_11),
    .io_wgt_data_bits_2_12(mvc_io_wgt_data_bits_2_12),
    .io_wgt_data_bits_2_13(mvc_io_wgt_data_bits_2_13),
    .io_wgt_data_bits_2_14(mvc_io_wgt_data_bits_2_14),
    .io_wgt_data_bits_2_15(mvc_io_wgt_data_bits_2_15),
    .io_wgt_data_bits_3_0(mvc_io_wgt_data_bits_3_0),
    .io_wgt_data_bits_3_1(mvc_io_wgt_data_bits_3_1),
    .io_wgt_data_bits_3_2(mvc_io_wgt_data_bits_3_2),
    .io_wgt_data_bits_3_3(mvc_io_wgt_data_bits_3_3),
    .io_wgt_data_bits_3_4(mvc_io_wgt_data_bits_3_4),
    .io_wgt_data_bits_3_5(mvc_io_wgt_data_bits_3_5),
    .io_wgt_data_bits_3_6(mvc_io_wgt_data_bits_3_6),
    .io_wgt_data_bits_3_7(mvc_io_wgt_data_bits_3_7),
    .io_wgt_data_bits_3_8(mvc_io_wgt_data_bits_3_8),
    .io_wgt_data_bits_3_9(mvc_io_wgt_data_bits_3_9),
    .io_wgt_data_bits_3_10(mvc_io_wgt_data_bits_3_10),
    .io_wgt_data_bits_3_11(mvc_io_wgt_data_bits_3_11),
    .io_wgt_data_bits_3_12(mvc_io_wgt_data_bits_3_12),
    .io_wgt_data_bits_3_13(mvc_io_wgt_data_bits_3_13),
    .io_wgt_data_bits_3_14(mvc_io_wgt_data_bits_3_14),
    .io_wgt_data_bits_3_15(mvc_io_wgt_data_bits_3_15),
    .io_wgt_data_bits_4_0(mvc_io_wgt_data_bits_4_0),
    .io_wgt_data_bits_4_1(mvc_io_wgt_data_bits_4_1),
    .io_wgt_data_bits_4_2(mvc_io_wgt_data_bits_4_2),
    .io_wgt_data_bits_4_3(mvc_io_wgt_data_bits_4_3),
    .io_wgt_data_bits_4_4(mvc_io_wgt_data_bits_4_4),
    .io_wgt_data_bits_4_5(mvc_io_wgt_data_bits_4_5),
    .io_wgt_data_bits_4_6(mvc_io_wgt_data_bits_4_6),
    .io_wgt_data_bits_4_7(mvc_io_wgt_data_bits_4_7),
    .io_wgt_data_bits_4_8(mvc_io_wgt_data_bits_4_8),
    .io_wgt_data_bits_4_9(mvc_io_wgt_data_bits_4_9),
    .io_wgt_data_bits_4_10(mvc_io_wgt_data_bits_4_10),
    .io_wgt_data_bits_4_11(mvc_io_wgt_data_bits_4_11),
    .io_wgt_data_bits_4_12(mvc_io_wgt_data_bits_4_12),
    .io_wgt_data_bits_4_13(mvc_io_wgt_data_bits_4_13),
    .io_wgt_data_bits_4_14(mvc_io_wgt_data_bits_4_14),
    .io_wgt_data_bits_4_15(mvc_io_wgt_data_bits_4_15),
    .io_wgt_data_bits_5_0(mvc_io_wgt_data_bits_5_0),
    .io_wgt_data_bits_5_1(mvc_io_wgt_data_bits_5_1),
    .io_wgt_data_bits_5_2(mvc_io_wgt_data_bits_5_2),
    .io_wgt_data_bits_5_3(mvc_io_wgt_data_bits_5_3),
    .io_wgt_data_bits_5_4(mvc_io_wgt_data_bits_5_4),
    .io_wgt_data_bits_5_5(mvc_io_wgt_data_bits_5_5),
    .io_wgt_data_bits_5_6(mvc_io_wgt_data_bits_5_6),
    .io_wgt_data_bits_5_7(mvc_io_wgt_data_bits_5_7),
    .io_wgt_data_bits_5_8(mvc_io_wgt_data_bits_5_8),
    .io_wgt_data_bits_5_9(mvc_io_wgt_data_bits_5_9),
    .io_wgt_data_bits_5_10(mvc_io_wgt_data_bits_5_10),
    .io_wgt_data_bits_5_11(mvc_io_wgt_data_bits_5_11),
    .io_wgt_data_bits_5_12(mvc_io_wgt_data_bits_5_12),
    .io_wgt_data_bits_5_13(mvc_io_wgt_data_bits_5_13),
    .io_wgt_data_bits_5_14(mvc_io_wgt_data_bits_5_14),
    .io_wgt_data_bits_5_15(mvc_io_wgt_data_bits_5_15),
    .io_wgt_data_bits_6_0(mvc_io_wgt_data_bits_6_0),
    .io_wgt_data_bits_6_1(mvc_io_wgt_data_bits_6_1),
    .io_wgt_data_bits_6_2(mvc_io_wgt_data_bits_6_2),
    .io_wgt_data_bits_6_3(mvc_io_wgt_data_bits_6_3),
    .io_wgt_data_bits_6_4(mvc_io_wgt_data_bits_6_4),
    .io_wgt_data_bits_6_5(mvc_io_wgt_data_bits_6_5),
    .io_wgt_data_bits_6_6(mvc_io_wgt_data_bits_6_6),
    .io_wgt_data_bits_6_7(mvc_io_wgt_data_bits_6_7),
    .io_wgt_data_bits_6_8(mvc_io_wgt_data_bits_6_8),
    .io_wgt_data_bits_6_9(mvc_io_wgt_data_bits_6_9),
    .io_wgt_data_bits_6_10(mvc_io_wgt_data_bits_6_10),
    .io_wgt_data_bits_6_11(mvc_io_wgt_data_bits_6_11),
    .io_wgt_data_bits_6_12(mvc_io_wgt_data_bits_6_12),
    .io_wgt_data_bits_6_13(mvc_io_wgt_data_bits_6_13),
    .io_wgt_data_bits_6_14(mvc_io_wgt_data_bits_6_14),
    .io_wgt_data_bits_6_15(mvc_io_wgt_data_bits_6_15),
    .io_wgt_data_bits_7_0(mvc_io_wgt_data_bits_7_0),
    .io_wgt_data_bits_7_1(mvc_io_wgt_data_bits_7_1),
    .io_wgt_data_bits_7_2(mvc_io_wgt_data_bits_7_2),
    .io_wgt_data_bits_7_3(mvc_io_wgt_data_bits_7_3),
    .io_wgt_data_bits_7_4(mvc_io_wgt_data_bits_7_4),
    .io_wgt_data_bits_7_5(mvc_io_wgt_data_bits_7_5),
    .io_wgt_data_bits_7_6(mvc_io_wgt_data_bits_7_6),
    .io_wgt_data_bits_7_7(mvc_io_wgt_data_bits_7_7),
    .io_wgt_data_bits_7_8(mvc_io_wgt_data_bits_7_8),
    .io_wgt_data_bits_7_9(mvc_io_wgt_data_bits_7_9),
    .io_wgt_data_bits_7_10(mvc_io_wgt_data_bits_7_10),
    .io_wgt_data_bits_7_11(mvc_io_wgt_data_bits_7_11),
    .io_wgt_data_bits_7_12(mvc_io_wgt_data_bits_7_12),
    .io_wgt_data_bits_7_13(mvc_io_wgt_data_bits_7_13),
    .io_wgt_data_bits_7_14(mvc_io_wgt_data_bits_7_14),
    .io_wgt_data_bits_7_15(mvc_io_wgt_data_bits_7_15),
    .io_wgt_data_bits_8_0(mvc_io_wgt_data_bits_8_0),
    .io_wgt_data_bits_8_1(mvc_io_wgt_data_bits_8_1),
    .io_wgt_data_bits_8_2(mvc_io_wgt_data_bits_8_2),
    .io_wgt_data_bits_8_3(mvc_io_wgt_data_bits_8_3),
    .io_wgt_data_bits_8_4(mvc_io_wgt_data_bits_8_4),
    .io_wgt_data_bits_8_5(mvc_io_wgt_data_bits_8_5),
    .io_wgt_data_bits_8_6(mvc_io_wgt_data_bits_8_6),
    .io_wgt_data_bits_8_7(mvc_io_wgt_data_bits_8_7),
    .io_wgt_data_bits_8_8(mvc_io_wgt_data_bits_8_8),
    .io_wgt_data_bits_8_9(mvc_io_wgt_data_bits_8_9),
    .io_wgt_data_bits_8_10(mvc_io_wgt_data_bits_8_10),
    .io_wgt_data_bits_8_11(mvc_io_wgt_data_bits_8_11),
    .io_wgt_data_bits_8_12(mvc_io_wgt_data_bits_8_12),
    .io_wgt_data_bits_8_13(mvc_io_wgt_data_bits_8_13),
    .io_wgt_data_bits_8_14(mvc_io_wgt_data_bits_8_14),
    .io_wgt_data_bits_8_15(mvc_io_wgt_data_bits_8_15),
    .io_wgt_data_bits_9_0(mvc_io_wgt_data_bits_9_0),
    .io_wgt_data_bits_9_1(mvc_io_wgt_data_bits_9_1),
    .io_wgt_data_bits_9_2(mvc_io_wgt_data_bits_9_2),
    .io_wgt_data_bits_9_3(mvc_io_wgt_data_bits_9_3),
    .io_wgt_data_bits_9_4(mvc_io_wgt_data_bits_9_4),
    .io_wgt_data_bits_9_5(mvc_io_wgt_data_bits_9_5),
    .io_wgt_data_bits_9_6(mvc_io_wgt_data_bits_9_6),
    .io_wgt_data_bits_9_7(mvc_io_wgt_data_bits_9_7),
    .io_wgt_data_bits_9_8(mvc_io_wgt_data_bits_9_8),
    .io_wgt_data_bits_9_9(mvc_io_wgt_data_bits_9_9),
    .io_wgt_data_bits_9_10(mvc_io_wgt_data_bits_9_10),
    .io_wgt_data_bits_9_11(mvc_io_wgt_data_bits_9_11),
    .io_wgt_data_bits_9_12(mvc_io_wgt_data_bits_9_12),
    .io_wgt_data_bits_9_13(mvc_io_wgt_data_bits_9_13),
    .io_wgt_data_bits_9_14(mvc_io_wgt_data_bits_9_14),
    .io_wgt_data_bits_9_15(mvc_io_wgt_data_bits_9_15),
    .io_wgt_data_bits_10_0(mvc_io_wgt_data_bits_10_0),
    .io_wgt_data_bits_10_1(mvc_io_wgt_data_bits_10_1),
    .io_wgt_data_bits_10_2(mvc_io_wgt_data_bits_10_2),
    .io_wgt_data_bits_10_3(mvc_io_wgt_data_bits_10_3),
    .io_wgt_data_bits_10_4(mvc_io_wgt_data_bits_10_4),
    .io_wgt_data_bits_10_5(mvc_io_wgt_data_bits_10_5),
    .io_wgt_data_bits_10_6(mvc_io_wgt_data_bits_10_6),
    .io_wgt_data_bits_10_7(mvc_io_wgt_data_bits_10_7),
    .io_wgt_data_bits_10_8(mvc_io_wgt_data_bits_10_8),
    .io_wgt_data_bits_10_9(mvc_io_wgt_data_bits_10_9),
    .io_wgt_data_bits_10_10(mvc_io_wgt_data_bits_10_10),
    .io_wgt_data_bits_10_11(mvc_io_wgt_data_bits_10_11),
    .io_wgt_data_bits_10_12(mvc_io_wgt_data_bits_10_12),
    .io_wgt_data_bits_10_13(mvc_io_wgt_data_bits_10_13),
    .io_wgt_data_bits_10_14(mvc_io_wgt_data_bits_10_14),
    .io_wgt_data_bits_10_15(mvc_io_wgt_data_bits_10_15),
    .io_wgt_data_bits_11_0(mvc_io_wgt_data_bits_11_0),
    .io_wgt_data_bits_11_1(mvc_io_wgt_data_bits_11_1),
    .io_wgt_data_bits_11_2(mvc_io_wgt_data_bits_11_2),
    .io_wgt_data_bits_11_3(mvc_io_wgt_data_bits_11_3),
    .io_wgt_data_bits_11_4(mvc_io_wgt_data_bits_11_4),
    .io_wgt_data_bits_11_5(mvc_io_wgt_data_bits_11_5),
    .io_wgt_data_bits_11_6(mvc_io_wgt_data_bits_11_6),
    .io_wgt_data_bits_11_7(mvc_io_wgt_data_bits_11_7),
    .io_wgt_data_bits_11_8(mvc_io_wgt_data_bits_11_8),
    .io_wgt_data_bits_11_9(mvc_io_wgt_data_bits_11_9),
    .io_wgt_data_bits_11_10(mvc_io_wgt_data_bits_11_10),
    .io_wgt_data_bits_11_11(mvc_io_wgt_data_bits_11_11),
    .io_wgt_data_bits_11_12(mvc_io_wgt_data_bits_11_12),
    .io_wgt_data_bits_11_13(mvc_io_wgt_data_bits_11_13),
    .io_wgt_data_bits_11_14(mvc_io_wgt_data_bits_11_14),
    .io_wgt_data_bits_11_15(mvc_io_wgt_data_bits_11_15),
    .io_wgt_data_bits_12_0(mvc_io_wgt_data_bits_12_0),
    .io_wgt_data_bits_12_1(mvc_io_wgt_data_bits_12_1),
    .io_wgt_data_bits_12_2(mvc_io_wgt_data_bits_12_2),
    .io_wgt_data_bits_12_3(mvc_io_wgt_data_bits_12_3),
    .io_wgt_data_bits_12_4(mvc_io_wgt_data_bits_12_4),
    .io_wgt_data_bits_12_5(mvc_io_wgt_data_bits_12_5),
    .io_wgt_data_bits_12_6(mvc_io_wgt_data_bits_12_6),
    .io_wgt_data_bits_12_7(mvc_io_wgt_data_bits_12_7),
    .io_wgt_data_bits_12_8(mvc_io_wgt_data_bits_12_8),
    .io_wgt_data_bits_12_9(mvc_io_wgt_data_bits_12_9),
    .io_wgt_data_bits_12_10(mvc_io_wgt_data_bits_12_10),
    .io_wgt_data_bits_12_11(mvc_io_wgt_data_bits_12_11),
    .io_wgt_data_bits_12_12(mvc_io_wgt_data_bits_12_12),
    .io_wgt_data_bits_12_13(mvc_io_wgt_data_bits_12_13),
    .io_wgt_data_bits_12_14(mvc_io_wgt_data_bits_12_14),
    .io_wgt_data_bits_12_15(mvc_io_wgt_data_bits_12_15),
    .io_wgt_data_bits_13_0(mvc_io_wgt_data_bits_13_0),
    .io_wgt_data_bits_13_1(mvc_io_wgt_data_bits_13_1),
    .io_wgt_data_bits_13_2(mvc_io_wgt_data_bits_13_2),
    .io_wgt_data_bits_13_3(mvc_io_wgt_data_bits_13_3),
    .io_wgt_data_bits_13_4(mvc_io_wgt_data_bits_13_4),
    .io_wgt_data_bits_13_5(mvc_io_wgt_data_bits_13_5),
    .io_wgt_data_bits_13_6(mvc_io_wgt_data_bits_13_6),
    .io_wgt_data_bits_13_7(mvc_io_wgt_data_bits_13_7),
    .io_wgt_data_bits_13_8(mvc_io_wgt_data_bits_13_8),
    .io_wgt_data_bits_13_9(mvc_io_wgt_data_bits_13_9),
    .io_wgt_data_bits_13_10(mvc_io_wgt_data_bits_13_10),
    .io_wgt_data_bits_13_11(mvc_io_wgt_data_bits_13_11),
    .io_wgt_data_bits_13_12(mvc_io_wgt_data_bits_13_12),
    .io_wgt_data_bits_13_13(mvc_io_wgt_data_bits_13_13),
    .io_wgt_data_bits_13_14(mvc_io_wgt_data_bits_13_14),
    .io_wgt_data_bits_13_15(mvc_io_wgt_data_bits_13_15),
    .io_wgt_data_bits_14_0(mvc_io_wgt_data_bits_14_0),
    .io_wgt_data_bits_14_1(mvc_io_wgt_data_bits_14_1),
    .io_wgt_data_bits_14_2(mvc_io_wgt_data_bits_14_2),
    .io_wgt_data_bits_14_3(mvc_io_wgt_data_bits_14_3),
    .io_wgt_data_bits_14_4(mvc_io_wgt_data_bits_14_4),
    .io_wgt_data_bits_14_5(mvc_io_wgt_data_bits_14_5),
    .io_wgt_data_bits_14_6(mvc_io_wgt_data_bits_14_6),
    .io_wgt_data_bits_14_7(mvc_io_wgt_data_bits_14_7),
    .io_wgt_data_bits_14_8(mvc_io_wgt_data_bits_14_8),
    .io_wgt_data_bits_14_9(mvc_io_wgt_data_bits_14_9),
    .io_wgt_data_bits_14_10(mvc_io_wgt_data_bits_14_10),
    .io_wgt_data_bits_14_11(mvc_io_wgt_data_bits_14_11),
    .io_wgt_data_bits_14_12(mvc_io_wgt_data_bits_14_12),
    .io_wgt_data_bits_14_13(mvc_io_wgt_data_bits_14_13),
    .io_wgt_data_bits_14_14(mvc_io_wgt_data_bits_14_14),
    .io_wgt_data_bits_14_15(mvc_io_wgt_data_bits_14_15),
    .io_wgt_data_bits_15_0(mvc_io_wgt_data_bits_15_0),
    .io_wgt_data_bits_15_1(mvc_io_wgt_data_bits_15_1),
    .io_wgt_data_bits_15_2(mvc_io_wgt_data_bits_15_2),
    .io_wgt_data_bits_15_3(mvc_io_wgt_data_bits_15_3),
    .io_wgt_data_bits_15_4(mvc_io_wgt_data_bits_15_4),
    .io_wgt_data_bits_15_5(mvc_io_wgt_data_bits_15_5),
    .io_wgt_data_bits_15_6(mvc_io_wgt_data_bits_15_6),
    .io_wgt_data_bits_15_7(mvc_io_wgt_data_bits_15_7),
    .io_wgt_data_bits_15_8(mvc_io_wgt_data_bits_15_8),
    .io_wgt_data_bits_15_9(mvc_io_wgt_data_bits_15_9),
    .io_wgt_data_bits_15_10(mvc_io_wgt_data_bits_15_10),
    .io_wgt_data_bits_15_11(mvc_io_wgt_data_bits_15_11),
    .io_wgt_data_bits_15_12(mvc_io_wgt_data_bits_15_12),
    .io_wgt_data_bits_15_13(mvc_io_wgt_data_bits_15_13),
    .io_wgt_data_bits_15_14(mvc_io_wgt_data_bits_15_14),
    .io_wgt_data_bits_15_15(mvc_io_wgt_data_bits_15_15),
    .io_acc_i_data_valid(mvc_io_acc_i_data_valid),
    .io_acc_i_data_bits_0_0(mvc_io_acc_i_data_bits_0_0),
    .io_acc_i_data_bits_0_1(mvc_io_acc_i_data_bits_0_1),
    .io_acc_i_data_bits_0_2(mvc_io_acc_i_data_bits_0_2),
    .io_acc_i_data_bits_0_3(mvc_io_acc_i_data_bits_0_3),
    .io_acc_i_data_bits_0_4(mvc_io_acc_i_data_bits_0_4),
    .io_acc_i_data_bits_0_5(mvc_io_acc_i_data_bits_0_5),
    .io_acc_i_data_bits_0_6(mvc_io_acc_i_data_bits_0_6),
    .io_acc_i_data_bits_0_7(mvc_io_acc_i_data_bits_0_7),
    .io_acc_i_data_bits_0_8(mvc_io_acc_i_data_bits_0_8),
    .io_acc_i_data_bits_0_9(mvc_io_acc_i_data_bits_0_9),
    .io_acc_i_data_bits_0_10(mvc_io_acc_i_data_bits_0_10),
    .io_acc_i_data_bits_0_11(mvc_io_acc_i_data_bits_0_11),
    .io_acc_i_data_bits_0_12(mvc_io_acc_i_data_bits_0_12),
    .io_acc_i_data_bits_0_13(mvc_io_acc_i_data_bits_0_13),
    .io_acc_i_data_bits_0_14(mvc_io_acc_i_data_bits_0_14),
    .io_acc_i_data_bits_0_15(mvc_io_acc_i_data_bits_0_15),
    .io_acc_o_data_valid(mvc_io_acc_o_data_valid),
    .io_acc_o_data_bits_0_0(mvc_io_acc_o_data_bits_0_0),
    .io_acc_o_data_bits_0_1(mvc_io_acc_o_data_bits_0_1),
    .io_acc_o_data_bits_0_2(mvc_io_acc_o_data_bits_0_2),
    .io_acc_o_data_bits_0_3(mvc_io_acc_o_data_bits_0_3),
    .io_acc_o_data_bits_0_4(mvc_io_acc_o_data_bits_0_4),
    .io_acc_o_data_bits_0_5(mvc_io_acc_o_data_bits_0_5),
    .io_acc_o_data_bits_0_6(mvc_io_acc_o_data_bits_0_6),
    .io_acc_o_data_bits_0_7(mvc_io_acc_o_data_bits_0_7),
    .io_acc_o_data_bits_0_8(mvc_io_acc_o_data_bits_0_8),
    .io_acc_o_data_bits_0_9(mvc_io_acc_o_data_bits_0_9),
    .io_acc_o_data_bits_0_10(mvc_io_acc_o_data_bits_0_10),
    .io_acc_o_data_bits_0_11(mvc_io_acc_o_data_bits_0_11),
    .io_acc_o_data_bits_0_12(mvc_io_acc_o_data_bits_0_12),
    .io_acc_o_data_bits_0_13(mvc_io_acc_o_data_bits_0_13),
    .io_acc_o_data_bits_0_14(mvc_io_acc_o_data_bits_0_14),
    .io_acc_o_data_bits_0_15(mvc_io_acc_o_data_bits_0_15),
    .io_out_data_valid(mvc_io_out_data_valid),
    .io_out_data_bits_0_0(mvc_io_out_data_bits_0_0),
    .io_out_data_bits_0_1(mvc_io_out_data_bits_0_1),
    .io_out_data_bits_0_2(mvc_io_out_data_bits_0_2),
    .io_out_data_bits_0_3(mvc_io_out_data_bits_0_3),
    .io_out_data_bits_0_4(mvc_io_out_data_bits_0_4),
    .io_out_data_bits_0_5(mvc_io_out_data_bits_0_5),
    .io_out_data_bits_0_6(mvc_io_out_data_bits_0_6),
    .io_out_data_bits_0_7(mvc_io_out_data_bits_0_7),
    .io_out_data_bits_0_8(mvc_io_out_data_bits_0_8),
    .io_out_data_bits_0_9(mvc_io_out_data_bits_0_9),
    .io_out_data_bits_0_10(mvc_io_out_data_bits_0_10),
    .io_out_data_bits_0_11(mvc_io_out_data_bits_0_11),
    .io_out_data_bits_0_12(mvc_io_out_data_bits_0_12),
    .io_out_data_bits_0_13(mvc_io_out_data_bits_0_13),
    .io_out_data_bits_0_14(mvc_io_out_data_bits_0_14),
    .io_out_data_bits_0_15(mvc_io_out_data_bits_0_15)
  );
  Pipe_16 wrpipe ( // @[TensorGemm.scala 218:22:@20644.4]
    .clock(wrpipe_clock),
    .reset(wrpipe_reset),
    .io_enq_valid(wrpipe_io_enq_valid),
    .io_enq_bits(wrpipe_io_enq_bits),
    .io_deq_valid(wrpipe_io_deq_valid),
    .io_deq_bits(wrpipe_io_deq_bits)
  );
  assign dec_reset = io_inst[7]; // @[TensorGemm.scala 200:29:@20607.4]
  assign dec_uop_begin = io_inst[20:8]; // @[TensorGemm.scala 200:29:@20609.4]
  assign dec_uop_end = io_inst[34:21]; // @[TensorGemm.scala 200:29:@20611.4]
  assign dec_lp_0 = io_inst[48:35]; // @[TensorGemm.scala 200:29:@20613.4]
  assign dec_lp_1 = io_inst[62:49]; // @[TensorGemm.scala 200:29:@20615.4]
  assign dec_acc_0 = io_inst[74:64]; // @[TensorGemm.scala 200:29:@20619.4]
  assign dec_acc_1 = io_inst[85:75]; // @[TensorGemm.scala 200:29:@20621.4]
  assign dec_inp_0 = io_inst[96:86]; // @[TensorGemm.scala 200:29:@20623.4]
  assign dec_inp_1 = io_inst[107:97]; // @[TensorGemm.scala 200:29:@20625.4]
  assign dec_wgt_0 = io_inst[117:108]; // @[TensorGemm.scala 200:29:@20627.4]
  assign dec_wgt_1 = io_inst[127:118]; // @[TensorGemm.scala 200:29:@20629.4]
  assign _T_7688 = inflight == 5'h0; // @[TensorGemm.scala 219:23:@20647.4]
  assign _T_7689 = state == 3'h4; // @[TensorGemm.scala 220:13:@20648.4]
  assign _T_7691 = dec_lp_0 - 14'h1; // @[TensorGemm.scala 221:26:@20649.4]
  assign _T_7692 = $unsigned(_T_7691); // @[TensorGemm.scala 221:26:@20650.4]
  assign _T_7693 = _T_7692[13:0]; // @[TensorGemm.scala 221:26:@20651.4]
  assign _T_7694 = cnt_o == _T_7693; // @[TensorGemm.scala 221:13:@20652.4]
  assign _T_7695 = _T_7689 & _T_7694; // @[TensorGemm.scala 220:22:@20653.4]
  assign _T_7697 = dec_lp_1 - 14'h1; // @[TensorGemm.scala 222:26:@20654.4]
  assign _T_7698 = $unsigned(_T_7697); // @[TensorGemm.scala 222:26:@20655.4]
  assign _T_7699 = _T_7698[13:0]; // @[TensorGemm.scala 222:26:@20656.4]
  assign _T_7700 = cnt_i == _T_7699; // @[TensorGemm.scala 222:13:@20657.4]
  assign _T_7701 = _T_7695 & _T_7700; // @[TensorGemm.scala 221:32:@20658.4]
  assign _T_7703 = dec_uop_end - 14'h1; // @[TensorGemm.scala 223:27:@20659.4]
  assign _T_7704 = $unsigned(_T_7703); // @[TensorGemm.scala 223:27:@20660.4]
  assign _T_7705 = _T_7704[13:0]; // @[TensorGemm.scala 223:27:@20661.4]
  assign _T_7706 = uop_idx == _T_7705; // @[TensorGemm.scala 223:15:@20662.4]
  assign _T_7707 = _T_7701 & _T_7706; // @[TensorGemm.scala 222:32:@20663.4]
  assign _T_7710 = _T_7707 & _T_7688; // @[TensorGemm.scala 223:33:@20665.4]
  assign _T_7711 = state == 3'h5; // @[TensorGemm.scala 225:13:@20666.4]
  assign _T_7712 = _T_7710 | _T_7711; // @[TensorGemm.scala 224:25:@20667.4]
  assign _T_7713 = 3'h0 == state; // @[Conditional.scala 37:30:@20669.4]
  assign _GEN_0 = io_start ? 3'h1 : state; // @[TensorGemm.scala 229:22:@20671.6]
  assign _T_7714 = 3'h1 == state; // @[Conditional.scala 37:30:@20676.6]
  assign _T_7715 = 3'h2 == state; // @[Conditional.scala 37:30:@20681.8]
  assign _T_7716 = 3'h3 == state; // @[Conditional.scala 37:30:@20686.10]
  assign _T_7717 = 3'h4 == state; // @[Conditional.scala 37:30:@20691.12]
  assign _T_7728 = _T_7694 & _T_7700; // @[TensorGemm.scala 244:36:@20701.14]
  assign _T_7734 = _T_7728 & _T_7706; // @[TensorGemm.scala 245:38:@20706.14]
  assign _T_7736 = inflight != 5'h0; // @[TensorGemm.scala 247:23:@20708.16]
  assign _GEN_1 = _T_7736 ? 3'h5 : 3'h0; // @[TensorGemm.scala 247:32:@20709.16]
  assign _GEN_2 = _T_7734 ? _GEN_1 : 3'h1; // @[TensorGemm.scala 246:40:@20707.14]
  assign _T_7737 = 3'h5 == state; // @[Conditional.scala 37:30:@20721.14]
  assign _GEN_3 = _T_7688 ? 3'h0 : state; // @[TensorGemm.scala 257:30:@20724.16]
  assign _GEN_4 = _T_7737 ? _GEN_3 : state; // @[Conditional.scala 39:67:@20722.14]
  assign _GEN_5 = _T_7717 ? _GEN_2 : _GEN_4; // @[Conditional.scala 39:67:@20692.12]
  assign _GEN_6 = _T_7716 ? 3'h4 : _GEN_5; // @[Conditional.scala 39:67:@20687.10]
  assign _GEN_7 = _T_7715 ? 3'h3 : _GEN_6; // @[Conditional.scala 39:67:@20682.8]
  assign _GEN_8 = _T_7714 ? 3'h2 : _GEN_7; // @[Conditional.scala 39:67:@20677.6]
  assign _GEN_9 = _T_7713 ? _GEN_0 : _GEN_8; // @[Conditional.scala 40:58:@20670.4]
  assign _T_7740 = state == 3'h0; // @[TensorGemm.scala 263:14:@20728.4]
  assign _T_7743 = dec_reset == 1'h0; // @[TensorGemm.scala 265:14:@20733.6]
  assign _T_7744 = state == 3'h3; // @[TensorGemm.scala 266:17:@20735.8]
  assign _T_7745 = _T_7744 & mvc_io_acc_o_data_valid; // @[TensorGemm.scala 266:34:@20736.8]
  assign _T_7748 = inflight + 5'h1; // @[TensorGemm.scala 269:28:@20743.12]
  assign _T_7749 = inflight + 5'h1; // @[TensorGemm.scala 269:28:@20744.12]
  assign _T_7751 = inflight - 5'h1; // @[TensorGemm.scala 271:28:@20749.14]
  assign _T_7752 = $unsigned(_T_7751); // @[TensorGemm.scala 271:28:@20750.14]
  assign _T_7753 = _T_7752[4:0]; // @[TensorGemm.scala 271:28:@20751.14]
  assign _GEN_10 = mvc_io_acc_o_data_valid ? _T_7753 : inflight; // @[TensorGemm.scala 270:41:@20748.12]
  assign _GEN_11 = _T_7744 ? _T_7749 : _GEN_10; // @[TensorGemm.scala 268:39:@20742.10]
  assign _GEN_12 = _T_7745 ? inflight : _GEN_11; // @[TensorGemm.scala 266:62:@20737.8]
  assign _GEN_13 = _T_7743 ? _GEN_12 : inflight; // @[TensorGemm.scala 265:26:@20734.6]
  assign _T_7761 = _T_7689 & _T_7706; // @[TensorGemm.scala 277:23:@20761.4]
  assign _T_7762 = _T_7740 | _T_7761; // @[TensorGemm.scala 276:21:@20762.4]
  assign _GEN_40 = {{1'd0}, dec_uop_begin}; // @[TensorGemm.scala 280:46:@20768.6]
  assign _T_7764 = _GEN_40 != dec_uop_end; // @[TensorGemm.scala 280:46:@20768.6]
  assign _T_7765 = _T_7689 & _T_7764; // @[TensorGemm.scala 280:29:@20769.6]
  assign _T_7767 = uop_idx + 14'h1; // @[TensorGemm.scala 281:24:@20771.8]
  assign _T_7768 = uop_idx + 14'h1; // @[TensorGemm.scala 281:24:@20772.8]
  assign _GEN_15 = _T_7765 ? _T_7768 : uop_idx; // @[TensorGemm.scala 280:59:@20770.6]
  assign _T_7786 = _T_7761 & _T_7700; // @[TensorGemm.scala 291:33:@20793.6]
  assign _T_7788 = cnt_o + 14'h1; // @[TensorGemm.scala 293:20:@20795.8]
  assign _T_7789 = cnt_o + 14'h1; // @[TensorGemm.scala 293:20:@20796.8]
  assign _GEN_41 = {{3'd0}, dec_acc_0}; // @[TensorGemm.scala 294:20:@20798.8]
  assign _T_7790 = acc_o + _GEN_41; // @[TensorGemm.scala 294:20:@20798.8]
  assign _T_7791 = acc_o + _GEN_41; // @[TensorGemm.scala 294:20:@20799.8]
  assign _GEN_42 = {{3'd0}, dec_inp_0}; // @[TensorGemm.scala 295:20:@20801.8]
  assign _T_7792 = inp_o + _GEN_42; // @[TensorGemm.scala 295:20:@20801.8]
  assign _T_7793 = inp_o + _GEN_42; // @[TensorGemm.scala 295:20:@20802.8]
  assign _GEN_43 = {{4'd0}, dec_wgt_0}; // @[TensorGemm.scala 296:20:@20804.8]
  assign _T_7794 = wgt_o + _GEN_43; // @[TensorGemm.scala 296:20:@20804.8]
  assign _T_7795 = wgt_o + _GEN_43; // @[TensorGemm.scala 296:20:@20805.8]
  assign _GEN_17 = _T_7786 ? _T_7789 : cnt_o; // @[TensorGemm.scala 292:33:@20794.6]
  assign _GEN_18 = _T_7786 ? _T_7791 : acc_o; // @[TensorGemm.scala 292:33:@20794.6]
  assign _GEN_19 = _T_7786 ? _T_7793 : inp_o; // @[TensorGemm.scala 292:33:@20794.6]
  assign _GEN_20 = _T_7786 ? _T_7795 : wgt_o; // @[TensorGemm.scala 292:33:@20794.6]
  assign _T_7801 = state == 3'h1; // @[TensorGemm.scala 304:20:@20816.6]
  assign _T_7802 = cnt_i == dec_lp_1; // @[TensorGemm.scala 304:42:@20817.6]
  assign _T_7803 = _T_7801 & _T_7802; // @[TensorGemm.scala 304:33:@20818.6]
  assign _T_7813 = cnt_i + 14'h1; // @[TensorGemm.scala 310:20:@20833.10]
  assign _T_7814 = cnt_i + 14'h1; // @[TensorGemm.scala 310:20:@20834.10]
  assign _GEN_44 = {{3'd0}, dec_acc_1}; // @[TensorGemm.scala 311:20:@20836.10]
  assign _T_7815 = acc_i + _GEN_44; // @[TensorGemm.scala 311:20:@20836.10]
  assign _T_7816 = acc_i + _GEN_44; // @[TensorGemm.scala 311:20:@20837.10]
  assign _GEN_45 = {{3'd0}, dec_inp_1}; // @[TensorGemm.scala 312:20:@20839.10]
  assign _T_7817 = inp_i + _GEN_45; // @[TensorGemm.scala 312:20:@20839.10]
  assign _T_7818 = inp_i + _GEN_45; // @[TensorGemm.scala 312:20:@20840.10]
  assign _GEN_46 = {{4'd0}, dec_wgt_1}; // @[TensorGemm.scala 313:20:@20842.10]
  assign _T_7819 = wgt_i + _GEN_46; // @[TensorGemm.scala 313:20:@20842.10]
  assign _T_7820 = wgt_i + _GEN_46; // @[TensorGemm.scala 313:20:@20843.10]
  assign _GEN_25 = _T_7761 ? _T_7814 : cnt_i; // @[TensorGemm.scala 309:59:@20832.8]
  assign _GEN_26 = _T_7761 ? _T_7816 : acc_i; // @[TensorGemm.scala 309:59:@20832.8]
  assign _GEN_27 = _T_7761 ? _T_7818 : inp_i; // @[TensorGemm.scala 309:59:@20832.8]
  assign _GEN_28 = _T_7761 ? _T_7820 : wgt_i; // @[TensorGemm.scala 309:59:@20832.8]
  assign _GEN_29 = _T_7803 ? 14'h0 : _GEN_25; // @[TensorGemm.scala 304:56:@20819.6]
  assign _GEN_30 = _T_7803 ? acc_o : _GEN_26; // @[TensorGemm.scala 304:56:@20819.6]
  assign _GEN_31 = _T_7803 ? inp_o : _GEN_27; // @[TensorGemm.scala 304:56:@20819.6]
  assign _GEN_32 = _T_7803 ? wgt_o : _GEN_28; // @[TensorGemm.scala 304:56:@20819.6]
  assign _T_7821 = state == 3'h2; // @[TensorGemm.scala 316:14:@20846.4]
  assign _T_7822 = _T_7821 & io_uop_data_valid; // @[TensorGemm.scala 316:30:@20847.4]
  assign _GEN_47 = {{3'd0}, io_uop_data_bits_u0}; // @[TensorGemm.scala 317:36:@20849.6]
  assign _T_7823 = _GEN_47 + acc_i; // @[TensorGemm.scala 317:36:@20849.6]
  assign _T_7824 = _GEN_47 + acc_i; // @[TensorGemm.scala 317:36:@20850.6]
  assign _GEN_48 = {{3'd0}, io_uop_data_bits_u1}; // @[TensorGemm.scala 318:36:@20852.6]
  assign _T_7825 = _GEN_48 + inp_i; // @[TensorGemm.scala 318:36:@20852.6]
  assign _T_7826 = _GEN_48 + inp_i; // @[TensorGemm.scala 318:36:@20853.6]
  assign _GEN_49 = {{4'd0}, io_uop_data_bits_u2}; // @[TensorGemm.scala 319:36:@20855.6]
  assign _T_7827 = _GEN_49 + wgt_i; // @[TensorGemm.scala 319:36:@20855.6]
  assign _T_7828 = _GEN_49 + wgt_i; // @[TensorGemm.scala 319:36:@20856.6]
  assign _T_7830 = ~ dec_reset; // @[TensorGemm.scala 322:43:@20860.4]
  assign _T_8115 = dec_reset ? 1'h1 : wrpipe_io_deq_valid; // @[TensorGemm.scala 351:8:@21446.4]
  assign _T_8117 = dec_reset ? uop_acc : wrpipe_io_deq_bits; // @[TensorGemm.scala 352:28:@21449.4]
  assign io_done = _T_7688 & _T_7712; // @[TensorGemm.scala 361:11:@21488.4]
  assign io_uop_idx_valid = state == 3'h1; // @[TensorGemm.scala 326:20:@20865.4]
  assign io_uop_idx_bits = uop_idx[10:0]; // @[TensorGemm.scala 327:19:@20866.4]
  assign io_inp_rd_idx_valid = state == 3'h3; // @[TensorGemm.scala 330:23:@20868.4]
  assign io_inp_rd_idx_bits = uop_inp[10:0]; // @[TensorGemm.scala 331:22:@20869.4]
  assign io_wgt_rd_idx_valid = state == 3'h3; // @[TensorGemm.scala 335:23:@20889.4]
  assign io_wgt_rd_idx_bits = uop_wgt[9:0]; // @[TensorGemm.scala 336:22:@20890.4]
  assign io_acc_rd_idx_valid = state == 3'h3; // @[TensorGemm.scala 340:23:@21150.4]
  assign io_acc_rd_idx_bits = uop_acc[10:0]; // @[TensorGemm.scala 341:22:@21151.4]
  assign io_acc_wr_valid = mvc_io_acc_o_data_valid & _T_8115; // @[TensorGemm.scala 350:19:@21448.4]
  assign io_acc_wr_bits_idx = _T_8117[10:0]; // @[TensorGemm.scala 352:22:@21450.4]
  assign io_acc_wr_bits_data_0_0 = mvc_io_acc_o_data_bits_0_0; // @[TensorGemm.scala 353:23:@21451.4]
  assign io_acc_wr_bits_data_0_1 = mvc_io_acc_o_data_bits_0_1; // @[TensorGemm.scala 353:23:@21452.4]
  assign io_acc_wr_bits_data_0_2 = mvc_io_acc_o_data_bits_0_2; // @[TensorGemm.scala 353:23:@21453.4]
  assign io_acc_wr_bits_data_0_3 = mvc_io_acc_o_data_bits_0_3; // @[TensorGemm.scala 353:23:@21454.4]
  assign io_acc_wr_bits_data_0_4 = mvc_io_acc_o_data_bits_0_4; // @[TensorGemm.scala 353:23:@21455.4]
  assign io_acc_wr_bits_data_0_5 = mvc_io_acc_o_data_bits_0_5; // @[TensorGemm.scala 353:23:@21456.4]
  assign io_acc_wr_bits_data_0_6 = mvc_io_acc_o_data_bits_0_6; // @[TensorGemm.scala 353:23:@21457.4]
  assign io_acc_wr_bits_data_0_7 = mvc_io_acc_o_data_bits_0_7; // @[TensorGemm.scala 353:23:@21458.4]
  assign io_acc_wr_bits_data_0_8 = mvc_io_acc_o_data_bits_0_8; // @[TensorGemm.scala 353:23:@21459.4]
  assign io_acc_wr_bits_data_0_9 = mvc_io_acc_o_data_bits_0_9; // @[TensorGemm.scala 353:23:@21460.4]
  assign io_acc_wr_bits_data_0_10 = mvc_io_acc_o_data_bits_0_10; // @[TensorGemm.scala 353:23:@21461.4]
  assign io_acc_wr_bits_data_0_11 = mvc_io_acc_o_data_bits_0_11; // @[TensorGemm.scala 353:23:@21462.4]
  assign io_acc_wr_bits_data_0_12 = mvc_io_acc_o_data_bits_0_12; // @[TensorGemm.scala 353:23:@21463.4]
  assign io_acc_wr_bits_data_0_13 = mvc_io_acc_o_data_bits_0_13; // @[TensorGemm.scala 353:23:@21464.4]
  assign io_acc_wr_bits_data_0_14 = mvc_io_acc_o_data_bits_0_14; // @[TensorGemm.scala 353:23:@21465.4]
  assign io_acc_wr_bits_data_0_15 = mvc_io_acc_o_data_bits_0_15; // @[TensorGemm.scala 353:23:@21466.4]
  assign io_out_wr_valid = mvc_io_out_data_valid & wrpipe_io_deq_valid; // @[TensorGemm.scala 356:19:@21468.4]
  assign io_out_wr_bits_idx = wrpipe_io_deq_bits[10:0]; // @[TensorGemm.scala 357:22:@21469.4]
  assign io_out_wr_bits_data_0_0 = mvc_io_out_data_bits_0_0; // @[TensorGemm.scala 358:23:@21470.4]
  assign io_out_wr_bits_data_0_1 = mvc_io_out_data_bits_0_1; // @[TensorGemm.scala 358:23:@21471.4]
  assign io_out_wr_bits_data_0_2 = mvc_io_out_data_bits_0_2; // @[TensorGemm.scala 358:23:@21472.4]
  assign io_out_wr_bits_data_0_3 = mvc_io_out_data_bits_0_3; // @[TensorGemm.scala 358:23:@21473.4]
  assign io_out_wr_bits_data_0_4 = mvc_io_out_data_bits_0_4; // @[TensorGemm.scala 358:23:@21474.4]
  assign io_out_wr_bits_data_0_5 = mvc_io_out_data_bits_0_5; // @[TensorGemm.scala 358:23:@21475.4]
  assign io_out_wr_bits_data_0_6 = mvc_io_out_data_bits_0_6; // @[TensorGemm.scala 358:23:@21476.4]
  assign io_out_wr_bits_data_0_7 = mvc_io_out_data_bits_0_7; // @[TensorGemm.scala 358:23:@21477.4]
  assign io_out_wr_bits_data_0_8 = mvc_io_out_data_bits_0_8; // @[TensorGemm.scala 358:23:@21478.4]
  assign io_out_wr_bits_data_0_9 = mvc_io_out_data_bits_0_9; // @[TensorGemm.scala 358:23:@21479.4]
  assign io_out_wr_bits_data_0_10 = mvc_io_out_data_bits_0_10; // @[TensorGemm.scala 358:23:@21480.4]
  assign io_out_wr_bits_data_0_11 = mvc_io_out_data_bits_0_11; // @[TensorGemm.scala 358:23:@21481.4]
  assign io_out_wr_bits_data_0_12 = mvc_io_out_data_bits_0_12; // @[TensorGemm.scala 358:23:@21482.4]
  assign io_out_wr_bits_data_0_13 = mvc_io_out_data_bits_0_13; // @[TensorGemm.scala 358:23:@21483.4]
  assign io_out_wr_bits_data_0_14 = mvc_io_out_data_bits_0_14; // @[TensorGemm.scala 358:23:@21484.4]
  assign io_out_wr_bits_data_0_15 = mvc_io_out_data_bits_0_15; // @[TensorGemm.scala 358:23:@21485.4]
  assign mvc_clock = clock; // @[:@20592.4]
  assign mvc_reset = reset; // @[:@20593.4]
  assign mvc_io_reset = dec_reset & _T_7689; // @[TensorGemm.scala 344:16:@21154.4]
  assign mvc_io_inp_data_valid = io_inp_rd_data_valid; // @[TensorGemm.scala 345:19:@21171.4]
  assign mvc_io_inp_data_bits_0_0 = io_inp_rd_data_bits_0_0; // @[TensorGemm.scala 345:19:@21155.4]
  assign mvc_io_inp_data_bits_0_1 = io_inp_rd_data_bits_0_1; // @[TensorGemm.scala 345:19:@21156.4]
  assign mvc_io_inp_data_bits_0_2 = io_inp_rd_data_bits_0_2; // @[TensorGemm.scala 345:19:@21157.4]
  assign mvc_io_inp_data_bits_0_3 = io_inp_rd_data_bits_0_3; // @[TensorGemm.scala 345:19:@21158.4]
  assign mvc_io_inp_data_bits_0_4 = io_inp_rd_data_bits_0_4; // @[TensorGemm.scala 345:19:@21159.4]
  assign mvc_io_inp_data_bits_0_5 = io_inp_rd_data_bits_0_5; // @[TensorGemm.scala 345:19:@21160.4]
  assign mvc_io_inp_data_bits_0_6 = io_inp_rd_data_bits_0_6; // @[TensorGemm.scala 345:19:@21161.4]
  assign mvc_io_inp_data_bits_0_7 = io_inp_rd_data_bits_0_7; // @[TensorGemm.scala 345:19:@21162.4]
  assign mvc_io_inp_data_bits_0_8 = io_inp_rd_data_bits_0_8; // @[TensorGemm.scala 345:19:@21163.4]
  assign mvc_io_inp_data_bits_0_9 = io_inp_rd_data_bits_0_9; // @[TensorGemm.scala 345:19:@21164.4]
  assign mvc_io_inp_data_bits_0_10 = io_inp_rd_data_bits_0_10; // @[TensorGemm.scala 345:19:@21165.4]
  assign mvc_io_inp_data_bits_0_11 = io_inp_rd_data_bits_0_11; // @[TensorGemm.scala 345:19:@21166.4]
  assign mvc_io_inp_data_bits_0_12 = io_inp_rd_data_bits_0_12; // @[TensorGemm.scala 345:19:@21167.4]
  assign mvc_io_inp_data_bits_0_13 = io_inp_rd_data_bits_0_13; // @[TensorGemm.scala 345:19:@21168.4]
  assign mvc_io_inp_data_bits_0_14 = io_inp_rd_data_bits_0_14; // @[TensorGemm.scala 345:19:@21169.4]
  assign mvc_io_inp_data_bits_0_15 = io_inp_rd_data_bits_0_15; // @[TensorGemm.scala 345:19:@21170.4]
  assign mvc_io_wgt_data_valid = io_wgt_rd_data_valid; // @[TensorGemm.scala 346:19:@21428.4]
  assign mvc_io_wgt_data_bits_0_0 = io_wgt_rd_data_bits_0_0; // @[TensorGemm.scala 346:19:@21172.4]
  assign mvc_io_wgt_data_bits_0_1 = io_wgt_rd_data_bits_0_1; // @[TensorGemm.scala 346:19:@21173.4]
  assign mvc_io_wgt_data_bits_0_2 = io_wgt_rd_data_bits_0_2; // @[TensorGemm.scala 346:19:@21174.4]
  assign mvc_io_wgt_data_bits_0_3 = io_wgt_rd_data_bits_0_3; // @[TensorGemm.scala 346:19:@21175.4]
  assign mvc_io_wgt_data_bits_0_4 = io_wgt_rd_data_bits_0_4; // @[TensorGemm.scala 346:19:@21176.4]
  assign mvc_io_wgt_data_bits_0_5 = io_wgt_rd_data_bits_0_5; // @[TensorGemm.scala 346:19:@21177.4]
  assign mvc_io_wgt_data_bits_0_6 = io_wgt_rd_data_bits_0_6; // @[TensorGemm.scala 346:19:@21178.4]
  assign mvc_io_wgt_data_bits_0_7 = io_wgt_rd_data_bits_0_7; // @[TensorGemm.scala 346:19:@21179.4]
  assign mvc_io_wgt_data_bits_0_8 = io_wgt_rd_data_bits_0_8; // @[TensorGemm.scala 346:19:@21180.4]
  assign mvc_io_wgt_data_bits_0_9 = io_wgt_rd_data_bits_0_9; // @[TensorGemm.scala 346:19:@21181.4]
  assign mvc_io_wgt_data_bits_0_10 = io_wgt_rd_data_bits_0_10; // @[TensorGemm.scala 346:19:@21182.4]
  assign mvc_io_wgt_data_bits_0_11 = io_wgt_rd_data_bits_0_11; // @[TensorGemm.scala 346:19:@21183.4]
  assign mvc_io_wgt_data_bits_0_12 = io_wgt_rd_data_bits_0_12; // @[TensorGemm.scala 346:19:@21184.4]
  assign mvc_io_wgt_data_bits_0_13 = io_wgt_rd_data_bits_0_13; // @[TensorGemm.scala 346:19:@21185.4]
  assign mvc_io_wgt_data_bits_0_14 = io_wgt_rd_data_bits_0_14; // @[TensorGemm.scala 346:19:@21186.4]
  assign mvc_io_wgt_data_bits_0_15 = io_wgt_rd_data_bits_0_15; // @[TensorGemm.scala 346:19:@21187.4]
  assign mvc_io_wgt_data_bits_1_0 = io_wgt_rd_data_bits_1_0; // @[TensorGemm.scala 346:19:@21188.4]
  assign mvc_io_wgt_data_bits_1_1 = io_wgt_rd_data_bits_1_1; // @[TensorGemm.scala 346:19:@21189.4]
  assign mvc_io_wgt_data_bits_1_2 = io_wgt_rd_data_bits_1_2; // @[TensorGemm.scala 346:19:@21190.4]
  assign mvc_io_wgt_data_bits_1_3 = io_wgt_rd_data_bits_1_3; // @[TensorGemm.scala 346:19:@21191.4]
  assign mvc_io_wgt_data_bits_1_4 = io_wgt_rd_data_bits_1_4; // @[TensorGemm.scala 346:19:@21192.4]
  assign mvc_io_wgt_data_bits_1_5 = io_wgt_rd_data_bits_1_5; // @[TensorGemm.scala 346:19:@21193.4]
  assign mvc_io_wgt_data_bits_1_6 = io_wgt_rd_data_bits_1_6; // @[TensorGemm.scala 346:19:@21194.4]
  assign mvc_io_wgt_data_bits_1_7 = io_wgt_rd_data_bits_1_7; // @[TensorGemm.scala 346:19:@21195.4]
  assign mvc_io_wgt_data_bits_1_8 = io_wgt_rd_data_bits_1_8; // @[TensorGemm.scala 346:19:@21196.4]
  assign mvc_io_wgt_data_bits_1_9 = io_wgt_rd_data_bits_1_9; // @[TensorGemm.scala 346:19:@21197.4]
  assign mvc_io_wgt_data_bits_1_10 = io_wgt_rd_data_bits_1_10; // @[TensorGemm.scala 346:19:@21198.4]
  assign mvc_io_wgt_data_bits_1_11 = io_wgt_rd_data_bits_1_11; // @[TensorGemm.scala 346:19:@21199.4]
  assign mvc_io_wgt_data_bits_1_12 = io_wgt_rd_data_bits_1_12; // @[TensorGemm.scala 346:19:@21200.4]
  assign mvc_io_wgt_data_bits_1_13 = io_wgt_rd_data_bits_1_13; // @[TensorGemm.scala 346:19:@21201.4]
  assign mvc_io_wgt_data_bits_1_14 = io_wgt_rd_data_bits_1_14; // @[TensorGemm.scala 346:19:@21202.4]
  assign mvc_io_wgt_data_bits_1_15 = io_wgt_rd_data_bits_1_15; // @[TensorGemm.scala 346:19:@21203.4]
  assign mvc_io_wgt_data_bits_2_0 = io_wgt_rd_data_bits_2_0; // @[TensorGemm.scala 346:19:@21204.4]
  assign mvc_io_wgt_data_bits_2_1 = io_wgt_rd_data_bits_2_1; // @[TensorGemm.scala 346:19:@21205.4]
  assign mvc_io_wgt_data_bits_2_2 = io_wgt_rd_data_bits_2_2; // @[TensorGemm.scala 346:19:@21206.4]
  assign mvc_io_wgt_data_bits_2_3 = io_wgt_rd_data_bits_2_3; // @[TensorGemm.scala 346:19:@21207.4]
  assign mvc_io_wgt_data_bits_2_4 = io_wgt_rd_data_bits_2_4; // @[TensorGemm.scala 346:19:@21208.4]
  assign mvc_io_wgt_data_bits_2_5 = io_wgt_rd_data_bits_2_5; // @[TensorGemm.scala 346:19:@21209.4]
  assign mvc_io_wgt_data_bits_2_6 = io_wgt_rd_data_bits_2_6; // @[TensorGemm.scala 346:19:@21210.4]
  assign mvc_io_wgt_data_bits_2_7 = io_wgt_rd_data_bits_2_7; // @[TensorGemm.scala 346:19:@21211.4]
  assign mvc_io_wgt_data_bits_2_8 = io_wgt_rd_data_bits_2_8; // @[TensorGemm.scala 346:19:@21212.4]
  assign mvc_io_wgt_data_bits_2_9 = io_wgt_rd_data_bits_2_9; // @[TensorGemm.scala 346:19:@21213.4]
  assign mvc_io_wgt_data_bits_2_10 = io_wgt_rd_data_bits_2_10; // @[TensorGemm.scala 346:19:@21214.4]
  assign mvc_io_wgt_data_bits_2_11 = io_wgt_rd_data_bits_2_11; // @[TensorGemm.scala 346:19:@21215.4]
  assign mvc_io_wgt_data_bits_2_12 = io_wgt_rd_data_bits_2_12; // @[TensorGemm.scala 346:19:@21216.4]
  assign mvc_io_wgt_data_bits_2_13 = io_wgt_rd_data_bits_2_13; // @[TensorGemm.scala 346:19:@21217.4]
  assign mvc_io_wgt_data_bits_2_14 = io_wgt_rd_data_bits_2_14; // @[TensorGemm.scala 346:19:@21218.4]
  assign mvc_io_wgt_data_bits_2_15 = io_wgt_rd_data_bits_2_15; // @[TensorGemm.scala 346:19:@21219.4]
  assign mvc_io_wgt_data_bits_3_0 = io_wgt_rd_data_bits_3_0; // @[TensorGemm.scala 346:19:@21220.4]
  assign mvc_io_wgt_data_bits_3_1 = io_wgt_rd_data_bits_3_1; // @[TensorGemm.scala 346:19:@21221.4]
  assign mvc_io_wgt_data_bits_3_2 = io_wgt_rd_data_bits_3_2; // @[TensorGemm.scala 346:19:@21222.4]
  assign mvc_io_wgt_data_bits_3_3 = io_wgt_rd_data_bits_3_3; // @[TensorGemm.scala 346:19:@21223.4]
  assign mvc_io_wgt_data_bits_3_4 = io_wgt_rd_data_bits_3_4; // @[TensorGemm.scala 346:19:@21224.4]
  assign mvc_io_wgt_data_bits_3_5 = io_wgt_rd_data_bits_3_5; // @[TensorGemm.scala 346:19:@21225.4]
  assign mvc_io_wgt_data_bits_3_6 = io_wgt_rd_data_bits_3_6; // @[TensorGemm.scala 346:19:@21226.4]
  assign mvc_io_wgt_data_bits_3_7 = io_wgt_rd_data_bits_3_7; // @[TensorGemm.scala 346:19:@21227.4]
  assign mvc_io_wgt_data_bits_3_8 = io_wgt_rd_data_bits_3_8; // @[TensorGemm.scala 346:19:@21228.4]
  assign mvc_io_wgt_data_bits_3_9 = io_wgt_rd_data_bits_3_9; // @[TensorGemm.scala 346:19:@21229.4]
  assign mvc_io_wgt_data_bits_3_10 = io_wgt_rd_data_bits_3_10; // @[TensorGemm.scala 346:19:@21230.4]
  assign mvc_io_wgt_data_bits_3_11 = io_wgt_rd_data_bits_3_11; // @[TensorGemm.scala 346:19:@21231.4]
  assign mvc_io_wgt_data_bits_3_12 = io_wgt_rd_data_bits_3_12; // @[TensorGemm.scala 346:19:@21232.4]
  assign mvc_io_wgt_data_bits_3_13 = io_wgt_rd_data_bits_3_13; // @[TensorGemm.scala 346:19:@21233.4]
  assign mvc_io_wgt_data_bits_3_14 = io_wgt_rd_data_bits_3_14; // @[TensorGemm.scala 346:19:@21234.4]
  assign mvc_io_wgt_data_bits_3_15 = io_wgt_rd_data_bits_3_15; // @[TensorGemm.scala 346:19:@21235.4]
  assign mvc_io_wgt_data_bits_4_0 = io_wgt_rd_data_bits_4_0; // @[TensorGemm.scala 346:19:@21236.4]
  assign mvc_io_wgt_data_bits_4_1 = io_wgt_rd_data_bits_4_1; // @[TensorGemm.scala 346:19:@21237.4]
  assign mvc_io_wgt_data_bits_4_2 = io_wgt_rd_data_bits_4_2; // @[TensorGemm.scala 346:19:@21238.4]
  assign mvc_io_wgt_data_bits_4_3 = io_wgt_rd_data_bits_4_3; // @[TensorGemm.scala 346:19:@21239.4]
  assign mvc_io_wgt_data_bits_4_4 = io_wgt_rd_data_bits_4_4; // @[TensorGemm.scala 346:19:@21240.4]
  assign mvc_io_wgt_data_bits_4_5 = io_wgt_rd_data_bits_4_5; // @[TensorGemm.scala 346:19:@21241.4]
  assign mvc_io_wgt_data_bits_4_6 = io_wgt_rd_data_bits_4_6; // @[TensorGemm.scala 346:19:@21242.4]
  assign mvc_io_wgt_data_bits_4_7 = io_wgt_rd_data_bits_4_7; // @[TensorGemm.scala 346:19:@21243.4]
  assign mvc_io_wgt_data_bits_4_8 = io_wgt_rd_data_bits_4_8; // @[TensorGemm.scala 346:19:@21244.4]
  assign mvc_io_wgt_data_bits_4_9 = io_wgt_rd_data_bits_4_9; // @[TensorGemm.scala 346:19:@21245.4]
  assign mvc_io_wgt_data_bits_4_10 = io_wgt_rd_data_bits_4_10; // @[TensorGemm.scala 346:19:@21246.4]
  assign mvc_io_wgt_data_bits_4_11 = io_wgt_rd_data_bits_4_11; // @[TensorGemm.scala 346:19:@21247.4]
  assign mvc_io_wgt_data_bits_4_12 = io_wgt_rd_data_bits_4_12; // @[TensorGemm.scala 346:19:@21248.4]
  assign mvc_io_wgt_data_bits_4_13 = io_wgt_rd_data_bits_4_13; // @[TensorGemm.scala 346:19:@21249.4]
  assign mvc_io_wgt_data_bits_4_14 = io_wgt_rd_data_bits_4_14; // @[TensorGemm.scala 346:19:@21250.4]
  assign mvc_io_wgt_data_bits_4_15 = io_wgt_rd_data_bits_4_15; // @[TensorGemm.scala 346:19:@21251.4]
  assign mvc_io_wgt_data_bits_5_0 = io_wgt_rd_data_bits_5_0; // @[TensorGemm.scala 346:19:@21252.4]
  assign mvc_io_wgt_data_bits_5_1 = io_wgt_rd_data_bits_5_1; // @[TensorGemm.scala 346:19:@21253.4]
  assign mvc_io_wgt_data_bits_5_2 = io_wgt_rd_data_bits_5_2; // @[TensorGemm.scala 346:19:@21254.4]
  assign mvc_io_wgt_data_bits_5_3 = io_wgt_rd_data_bits_5_3; // @[TensorGemm.scala 346:19:@21255.4]
  assign mvc_io_wgt_data_bits_5_4 = io_wgt_rd_data_bits_5_4; // @[TensorGemm.scala 346:19:@21256.4]
  assign mvc_io_wgt_data_bits_5_5 = io_wgt_rd_data_bits_5_5; // @[TensorGemm.scala 346:19:@21257.4]
  assign mvc_io_wgt_data_bits_5_6 = io_wgt_rd_data_bits_5_6; // @[TensorGemm.scala 346:19:@21258.4]
  assign mvc_io_wgt_data_bits_5_7 = io_wgt_rd_data_bits_5_7; // @[TensorGemm.scala 346:19:@21259.4]
  assign mvc_io_wgt_data_bits_5_8 = io_wgt_rd_data_bits_5_8; // @[TensorGemm.scala 346:19:@21260.4]
  assign mvc_io_wgt_data_bits_5_9 = io_wgt_rd_data_bits_5_9; // @[TensorGemm.scala 346:19:@21261.4]
  assign mvc_io_wgt_data_bits_5_10 = io_wgt_rd_data_bits_5_10; // @[TensorGemm.scala 346:19:@21262.4]
  assign mvc_io_wgt_data_bits_5_11 = io_wgt_rd_data_bits_5_11; // @[TensorGemm.scala 346:19:@21263.4]
  assign mvc_io_wgt_data_bits_5_12 = io_wgt_rd_data_bits_5_12; // @[TensorGemm.scala 346:19:@21264.4]
  assign mvc_io_wgt_data_bits_5_13 = io_wgt_rd_data_bits_5_13; // @[TensorGemm.scala 346:19:@21265.4]
  assign mvc_io_wgt_data_bits_5_14 = io_wgt_rd_data_bits_5_14; // @[TensorGemm.scala 346:19:@21266.4]
  assign mvc_io_wgt_data_bits_5_15 = io_wgt_rd_data_bits_5_15; // @[TensorGemm.scala 346:19:@21267.4]
  assign mvc_io_wgt_data_bits_6_0 = io_wgt_rd_data_bits_6_0; // @[TensorGemm.scala 346:19:@21268.4]
  assign mvc_io_wgt_data_bits_6_1 = io_wgt_rd_data_bits_6_1; // @[TensorGemm.scala 346:19:@21269.4]
  assign mvc_io_wgt_data_bits_6_2 = io_wgt_rd_data_bits_6_2; // @[TensorGemm.scala 346:19:@21270.4]
  assign mvc_io_wgt_data_bits_6_3 = io_wgt_rd_data_bits_6_3; // @[TensorGemm.scala 346:19:@21271.4]
  assign mvc_io_wgt_data_bits_6_4 = io_wgt_rd_data_bits_6_4; // @[TensorGemm.scala 346:19:@21272.4]
  assign mvc_io_wgt_data_bits_6_5 = io_wgt_rd_data_bits_6_5; // @[TensorGemm.scala 346:19:@21273.4]
  assign mvc_io_wgt_data_bits_6_6 = io_wgt_rd_data_bits_6_6; // @[TensorGemm.scala 346:19:@21274.4]
  assign mvc_io_wgt_data_bits_6_7 = io_wgt_rd_data_bits_6_7; // @[TensorGemm.scala 346:19:@21275.4]
  assign mvc_io_wgt_data_bits_6_8 = io_wgt_rd_data_bits_6_8; // @[TensorGemm.scala 346:19:@21276.4]
  assign mvc_io_wgt_data_bits_6_9 = io_wgt_rd_data_bits_6_9; // @[TensorGemm.scala 346:19:@21277.4]
  assign mvc_io_wgt_data_bits_6_10 = io_wgt_rd_data_bits_6_10; // @[TensorGemm.scala 346:19:@21278.4]
  assign mvc_io_wgt_data_bits_6_11 = io_wgt_rd_data_bits_6_11; // @[TensorGemm.scala 346:19:@21279.4]
  assign mvc_io_wgt_data_bits_6_12 = io_wgt_rd_data_bits_6_12; // @[TensorGemm.scala 346:19:@21280.4]
  assign mvc_io_wgt_data_bits_6_13 = io_wgt_rd_data_bits_6_13; // @[TensorGemm.scala 346:19:@21281.4]
  assign mvc_io_wgt_data_bits_6_14 = io_wgt_rd_data_bits_6_14; // @[TensorGemm.scala 346:19:@21282.4]
  assign mvc_io_wgt_data_bits_6_15 = io_wgt_rd_data_bits_6_15; // @[TensorGemm.scala 346:19:@21283.4]
  assign mvc_io_wgt_data_bits_7_0 = io_wgt_rd_data_bits_7_0; // @[TensorGemm.scala 346:19:@21284.4]
  assign mvc_io_wgt_data_bits_7_1 = io_wgt_rd_data_bits_7_1; // @[TensorGemm.scala 346:19:@21285.4]
  assign mvc_io_wgt_data_bits_7_2 = io_wgt_rd_data_bits_7_2; // @[TensorGemm.scala 346:19:@21286.4]
  assign mvc_io_wgt_data_bits_7_3 = io_wgt_rd_data_bits_7_3; // @[TensorGemm.scala 346:19:@21287.4]
  assign mvc_io_wgt_data_bits_7_4 = io_wgt_rd_data_bits_7_4; // @[TensorGemm.scala 346:19:@21288.4]
  assign mvc_io_wgt_data_bits_7_5 = io_wgt_rd_data_bits_7_5; // @[TensorGemm.scala 346:19:@21289.4]
  assign mvc_io_wgt_data_bits_7_6 = io_wgt_rd_data_bits_7_6; // @[TensorGemm.scala 346:19:@21290.4]
  assign mvc_io_wgt_data_bits_7_7 = io_wgt_rd_data_bits_7_7; // @[TensorGemm.scala 346:19:@21291.4]
  assign mvc_io_wgt_data_bits_7_8 = io_wgt_rd_data_bits_7_8; // @[TensorGemm.scala 346:19:@21292.4]
  assign mvc_io_wgt_data_bits_7_9 = io_wgt_rd_data_bits_7_9; // @[TensorGemm.scala 346:19:@21293.4]
  assign mvc_io_wgt_data_bits_7_10 = io_wgt_rd_data_bits_7_10; // @[TensorGemm.scala 346:19:@21294.4]
  assign mvc_io_wgt_data_bits_7_11 = io_wgt_rd_data_bits_7_11; // @[TensorGemm.scala 346:19:@21295.4]
  assign mvc_io_wgt_data_bits_7_12 = io_wgt_rd_data_bits_7_12; // @[TensorGemm.scala 346:19:@21296.4]
  assign mvc_io_wgt_data_bits_7_13 = io_wgt_rd_data_bits_7_13; // @[TensorGemm.scala 346:19:@21297.4]
  assign mvc_io_wgt_data_bits_7_14 = io_wgt_rd_data_bits_7_14; // @[TensorGemm.scala 346:19:@21298.4]
  assign mvc_io_wgt_data_bits_7_15 = io_wgt_rd_data_bits_7_15; // @[TensorGemm.scala 346:19:@21299.4]
  assign mvc_io_wgt_data_bits_8_0 = io_wgt_rd_data_bits_8_0; // @[TensorGemm.scala 346:19:@21300.4]
  assign mvc_io_wgt_data_bits_8_1 = io_wgt_rd_data_bits_8_1; // @[TensorGemm.scala 346:19:@21301.4]
  assign mvc_io_wgt_data_bits_8_2 = io_wgt_rd_data_bits_8_2; // @[TensorGemm.scala 346:19:@21302.4]
  assign mvc_io_wgt_data_bits_8_3 = io_wgt_rd_data_bits_8_3; // @[TensorGemm.scala 346:19:@21303.4]
  assign mvc_io_wgt_data_bits_8_4 = io_wgt_rd_data_bits_8_4; // @[TensorGemm.scala 346:19:@21304.4]
  assign mvc_io_wgt_data_bits_8_5 = io_wgt_rd_data_bits_8_5; // @[TensorGemm.scala 346:19:@21305.4]
  assign mvc_io_wgt_data_bits_8_6 = io_wgt_rd_data_bits_8_6; // @[TensorGemm.scala 346:19:@21306.4]
  assign mvc_io_wgt_data_bits_8_7 = io_wgt_rd_data_bits_8_7; // @[TensorGemm.scala 346:19:@21307.4]
  assign mvc_io_wgt_data_bits_8_8 = io_wgt_rd_data_bits_8_8; // @[TensorGemm.scala 346:19:@21308.4]
  assign mvc_io_wgt_data_bits_8_9 = io_wgt_rd_data_bits_8_9; // @[TensorGemm.scala 346:19:@21309.4]
  assign mvc_io_wgt_data_bits_8_10 = io_wgt_rd_data_bits_8_10; // @[TensorGemm.scala 346:19:@21310.4]
  assign mvc_io_wgt_data_bits_8_11 = io_wgt_rd_data_bits_8_11; // @[TensorGemm.scala 346:19:@21311.4]
  assign mvc_io_wgt_data_bits_8_12 = io_wgt_rd_data_bits_8_12; // @[TensorGemm.scala 346:19:@21312.4]
  assign mvc_io_wgt_data_bits_8_13 = io_wgt_rd_data_bits_8_13; // @[TensorGemm.scala 346:19:@21313.4]
  assign mvc_io_wgt_data_bits_8_14 = io_wgt_rd_data_bits_8_14; // @[TensorGemm.scala 346:19:@21314.4]
  assign mvc_io_wgt_data_bits_8_15 = io_wgt_rd_data_bits_8_15; // @[TensorGemm.scala 346:19:@21315.4]
  assign mvc_io_wgt_data_bits_9_0 = io_wgt_rd_data_bits_9_0; // @[TensorGemm.scala 346:19:@21316.4]
  assign mvc_io_wgt_data_bits_9_1 = io_wgt_rd_data_bits_9_1; // @[TensorGemm.scala 346:19:@21317.4]
  assign mvc_io_wgt_data_bits_9_2 = io_wgt_rd_data_bits_9_2; // @[TensorGemm.scala 346:19:@21318.4]
  assign mvc_io_wgt_data_bits_9_3 = io_wgt_rd_data_bits_9_3; // @[TensorGemm.scala 346:19:@21319.4]
  assign mvc_io_wgt_data_bits_9_4 = io_wgt_rd_data_bits_9_4; // @[TensorGemm.scala 346:19:@21320.4]
  assign mvc_io_wgt_data_bits_9_5 = io_wgt_rd_data_bits_9_5; // @[TensorGemm.scala 346:19:@21321.4]
  assign mvc_io_wgt_data_bits_9_6 = io_wgt_rd_data_bits_9_6; // @[TensorGemm.scala 346:19:@21322.4]
  assign mvc_io_wgt_data_bits_9_7 = io_wgt_rd_data_bits_9_7; // @[TensorGemm.scala 346:19:@21323.4]
  assign mvc_io_wgt_data_bits_9_8 = io_wgt_rd_data_bits_9_8; // @[TensorGemm.scala 346:19:@21324.4]
  assign mvc_io_wgt_data_bits_9_9 = io_wgt_rd_data_bits_9_9; // @[TensorGemm.scala 346:19:@21325.4]
  assign mvc_io_wgt_data_bits_9_10 = io_wgt_rd_data_bits_9_10; // @[TensorGemm.scala 346:19:@21326.4]
  assign mvc_io_wgt_data_bits_9_11 = io_wgt_rd_data_bits_9_11; // @[TensorGemm.scala 346:19:@21327.4]
  assign mvc_io_wgt_data_bits_9_12 = io_wgt_rd_data_bits_9_12; // @[TensorGemm.scala 346:19:@21328.4]
  assign mvc_io_wgt_data_bits_9_13 = io_wgt_rd_data_bits_9_13; // @[TensorGemm.scala 346:19:@21329.4]
  assign mvc_io_wgt_data_bits_9_14 = io_wgt_rd_data_bits_9_14; // @[TensorGemm.scala 346:19:@21330.4]
  assign mvc_io_wgt_data_bits_9_15 = io_wgt_rd_data_bits_9_15; // @[TensorGemm.scala 346:19:@21331.4]
  assign mvc_io_wgt_data_bits_10_0 = io_wgt_rd_data_bits_10_0; // @[TensorGemm.scala 346:19:@21332.4]
  assign mvc_io_wgt_data_bits_10_1 = io_wgt_rd_data_bits_10_1; // @[TensorGemm.scala 346:19:@21333.4]
  assign mvc_io_wgt_data_bits_10_2 = io_wgt_rd_data_bits_10_2; // @[TensorGemm.scala 346:19:@21334.4]
  assign mvc_io_wgt_data_bits_10_3 = io_wgt_rd_data_bits_10_3; // @[TensorGemm.scala 346:19:@21335.4]
  assign mvc_io_wgt_data_bits_10_4 = io_wgt_rd_data_bits_10_4; // @[TensorGemm.scala 346:19:@21336.4]
  assign mvc_io_wgt_data_bits_10_5 = io_wgt_rd_data_bits_10_5; // @[TensorGemm.scala 346:19:@21337.4]
  assign mvc_io_wgt_data_bits_10_6 = io_wgt_rd_data_bits_10_6; // @[TensorGemm.scala 346:19:@21338.4]
  assign mvc_io_wgt_data_bits_10_7 = io_wgt_rd_data_bits_10_7; // @[TensorGemm.scala 346:19:@21339.4]
  assign mvc_io_wgt_data_bits_10_8 = io_wgt_rd_data_bits_10_8; // @[TensorGemm.scala 346:19:@21340.4]
  assign mvc_io_wgt_data_bits_10_9 = io_wgt_rd_data_bits_10_9; // @[TensorGemm.scala 346:19:@21341.4]
  assign mvc_io_wgt_data_bits_10_10 = io_wgt_rd_data_bits_10_10; // @[TensorGemm.scala 346:19:@21342.4]
  assign mvc_io_wgt_data_bits_10_11 = io_wgt_rd_data_bits_10_11; // @[TensorGemm.scala 346:19:@21343.4]
  assign mvc_io_wgt_data_bits_10_12 = io_wgt_rd_data_bits_10_12; // @[TensorGemm.scala 346:19:@21344.4]
  assign mvc_io_wgt_data_bits_10_13 = io_wgt_rd_data_bits_10_13; // @[TensorGemm.scala 346:19:@21345.4]
  assign mvc_io_wgt_data_bits_10_14 = io_wgt_rd_data_bits_10_14; // @[TensorGemm.scala 346:19:@21346.4]
  assign mvc_io_wgt_data_bits_10_15 = io_wgt_rd_data_bits_10_15; // @[TensorGemm.scala 346:19:@21347.4]
  assign mvc_io_wgt_data_bits_11_0 = io_wgt_rd_data_bits_11_0; // @[TensorGemm.scala 346:19:@21348.4]
  assign mvc_io_wgt_data_bits_11_1 = io_wgt_rd_data_bits_11_1; // @[TensorGemm.scala 346:19:@21349.4]
  assign mvc_io_wgt_data_bits_11_2 = io_wgt_rd_data_bits_11_2; // @[TensorGemm.scala 346:19:@21350.4]
  assign mvc_io_wgt_data_bits_11_3 = io_wgt_rd_data_bits_11_3; // @[TensorGemm.scala 346:19:@21351.4]
  assign mvc_io_wgt_data_bits_11_4 = io_wgt_rd_data_bits_11_4; // @[TensorGemm.scala 346:19:@21352.4]
  assign mvc_io_wgt_data_bits_11_5 = io_wgt_rd_data_bits_11_5; // @[TensorGemm.scala 346:19:@21353.4]
  assign mvc_io_wgt_data_bits_11_6 = io_wgt_rd_data_bits_11_6; // @[TensorGemm.scala 346:19:@21354.4]
  assign mvc_io_wgt_data_bits_11_7 = io_wgt_rd_data_bits_11_7; // @[TensorGemm.scala 346:19:@21355.4]
  assign mvc_io_wgt_data_bits_11_8 = io_wgt_rd_data_bits_11_8; // @[TensorGemm.scala 346:19:@21356.4]
  assign mvc_io_wgt_data_bits_11_9 = io_wgt_rd_data_bits_11_9; // @[TensorGemm.scala 346:19:@21357.4]
  assign mvc_io_wgt_data_bits_11_10 = io_wgt_rd_data_bits_11_10; // @[TensorGemm.scala 346:19:@21358.4]
  assign mvc_io_wgt_data_bits_11_11 = io_wgt_rd_data_bits_11_11; // @[TensorGemm.scala 346:19:@21359.4]
  assign mvc_io_wgt_data_bits_11_12 = io_wgt_rd_data_bits_11_12; // @[TensorGemm.scala 346:19:@21360.4]
  assign mvc_io_wgt_data_bits_11_13 = io_wgt_rd_data_bits_11_13; // @[TensorGemm.scala 346:19:@21361.4]
  assign mvc_io_wgt_data_bits_11_14 = io_wgt_rd_data_bits_11_14; // @[TensorGemm.scala 346:19:@21362.4]
  assign mvc_io_wgt_data_bits_11_15 = io_wgt_rd_data_bits_11_15; // @[TensorGemm.scala 346:19:@21363.4]
  assign mvc_io_wgt_data_bits_12_0 = io_wgt_rd_data_bits_12_0; // @[TensorGemm.scala 346:19:@21364.4]
  assign mvc_io_wgt_data_bits_12_1 = io_wgt_rd_data_bits_12_1; // @[TensorGemm.scala 346:19:@21365.4]
  assign mvc_io_wgt_data_bits_12_2 = io_wgt_rd_data_bits_12_2; // @[TensorGemm.scala 346:19:@21366.4]
  assign mvc_io_wgt_data_bits_12_3 = io_wgt_rd_data_bits_12_3; // @[TensorGemm.scala 346:19:@21367.4]
  assign mvc_io_wgt_data_bits_12_4 = io_wgt_rd_data_bits_12_4; // @[TensorGemm.scala 346:19:@21368.4]
  assign mvc_io_wgt_data_bits_12_5 = io_wgt_rd_data_bits_12_5; // @[TensorGemm.scala 346:19:@21369.4]
  assign mvc_io_wgt_data_bits_12_6 = io_wgt_rd_data_bits_12_6; // @[TensorGemm.scala 346:19:@21370.4]
  assign mvc_io_wgt_data_bits_12_7 = io_wgt_rd_data_bits_12_7; // @[TensorGemm.scala 346:19:@21371.4]
  assign mvc_io_wgt_data_bits_12_8 = io_wgt_rd_data_bits_12_8; // @[TensorGemm.scala 346:19:@21372.4]
  assign mvc_io_wgt_data_bits_12_9 = io_wgt_rd_data_bits_12_9; // @[TensorGemm.scala 346:19:@21373.4]
  assign mvc_io_wgt_data_bits_12_10 = io_wgt_rd_data_bits_12_10; // @[TensorGemm.scala 346:19:@21374.4]
  assign mvc_io_wgt_data_bits_12_11 = io_wgt_rd_data_bits_12_11; // @[TensorGemm.scala 346:19:@21375.4]
  assign mvc_io_wgt_data_bits_12_12 = io_wgt_rd_data_bits_12_12; // @[TensorGemm.scala 346:19:@21376.4]
  assign mvc_io_wgt_data_bits_12_13 = io_wgt_rd_data_bits_12_13; // @[TensorGemm.scala 346:19:@21377.4]
  assign mvc_io_wgt_data_bits_12_14 = io_wgt_rd_data_bits_12_14; // @[TensorGemm.scala 346:19:@21378.4]
  assign mvc_io_wgt_data_bits_12_15 = io_wgt_rd_data_bits_12_15; // @[TensorGemm.scala 346:19:@21379.4]
  assign mvc_io_wgt_data_bits_13_0 = io_wgt_rd_data_bits_13_0; // @[TensorGemm.scala 346:19:@21380.4]
  assign mvc_io_wgt_data_bits_13_1 = io_wgt_rd_data_bits_13_1; // @[TensorGemm.scala 346:19:@21381.4]
  assign mvc_io_wgt_data_bits_13_2 = io_wgt_rd_data_bits_13_2; // @[TensorGemm.scala 346:19:@21382.4]
  assign mvc_io_wgt_data_bits_13_3 = io_wgt_rd_data_bits_13_3; // @[TensorGemm.scala 346:19:@21383.4]
  assign mvc_io_wgt_data_bits_13_4 = io_wgt_rd_data_bits_13_4; // @[TensorGemm.scala 346:19:@21384.4]
  assign mvc_io_wgt_data_bits_13_5 = io_wgt_rd_data_bits_13_5; // @[TensorGemm.scala 346:19:@21385.4]
  assign mvc_io_wgt_data_bits_13_6 = io_wgt_rd_data_bits_13_6; // @[TensorGemm.scala 346:19:@21386.4]
  assign mvc_io_wgt_data_bits_13_7 = io_wgt_rd_data_bits_13_7; // @[TensorGemm.scala 346:19:@21387.4]
  assign mvc_io_wgt_data_bits_13_8 = io_wgt_rd_data_bits_13_8; // @[TensorGemm.scala 346:19:@21388.4]
  assign mvc_io_wgt_data_bits_13_9 = io_wgt_rd_data_bits_13_9; // @[TensorGemm.scala 346:19:@21389.4]
  assign mvc_io_wgt_data_bits_13_10 = io_wgt_rd_data_bits_13_10; // @[TensorGemm.scala 346:19:@21390.4]
  assign mvc_io_wgt_data_bits_13_11 = io_wgt_rd_data_bits_13_11; // @[TensorGemm.scala 346:19:@21391.4]
  assign mvc_io_wgt_data_bits_13_12 = io_wgt_rd_data_bits_13_12; // @[TensorGemm.scala 346:19:@21392.4]
  assign mvc_io_wgt_data_bits_13_13 = io_wgt_rd_data_bits_13_13; // @[TensorGemm.scala 346:19:@21393.4]
  assign mvc_io_wgt_data_bits_13_14 = io_wgt_rd_data_bits_13_14; // @[TensorGemm.scala 346:19:@21394.4]
  assign mvc_io_wgt_data_bits_13_15 = io_wgt_rd_data_bits_13_15; // @[TensorGemm.scala 346:19:@21395.4]
  assign mvc_io_wgt_data_bits_14_0 = io_wgt_rd_data_bits_14_0; // @[TensorGemm.scala 346:19:@21396.4]
  assign mvc_io_wgt_data_bits_14_1 = io_wgt_rd_data_bits_14_1; // @[TensorGemm.scala 346:19:@21397.4]
  assign mvc_io_wgt_data_bits_14_2 = io_wgt_rd_data_bits_14_2; // @[TensorGemm.scala 346:19:@21398.4]
  assign mvc_io_wgt_data_bits_14_3 = io_wgt_rd_data_bits_14_3; // @[TensorGemm.scala 346:19:@21399.4]
  assign mvc_io_wgt_data_bits_14_4 = io_wgt_rd_data_bits_14_4; // @[TensorGemm.scala 346:19:@21400.4]
  assign mvc_io_wgt_data_bits_14_5 = io_wgt_rd_data_bits_14_5; // @[TensorGemm.scala 346:19:@21401.4]
  assign mvc_io_wgt_data_bits_14_6 = io_wgt_rd_data_bits_14_6; // @[TensorGemm.scala 346:19:@21402.4]
  assign mvc_io_wgt_data_bits_14_7 = io_wgt_rd_data_bits_14_7; // @[TensorGemm.scala 346:19:@21403.4]
  assign mvc_io_wgt_data_bits_14_8 = io_wgt_rd_data_bits_14_8; // @[TensorGemm.scala 346:19:@21404.4]
  assign mvc_io_wgt_data_bits_14_9 = io_wgt_rd_data_bits_14_9; // @[TensorGemm.scala 346:19:@21405.4]
  assign mvc_io_wgt_data_bits_14_10 = io_wgt_rd_data_bits_14_10; // @[TensorGemm.scala 346:19:@21406.4]
  assign mvc_io_wgt_data_bits_14_11 = io_wgt_rd_data_bits_14_11; // @[TensorGemm.scala 346:19:@21407.4]
  assign mvc_io_wgt_data_bits_14_12 = io_wgt_rd_data_bits_14_12; // @[TensorGemm.scala 346:19:@21408.4]
  assign mvc_io_wgt_data_bits_14_13 = io_wgt_rd_data_bits_14_13; // @[TensorGemm.scala 346:19:@21409.4]
  assign mvc_io_wgt_data_bits_14_14 = io_wgt_rd_data_bits_14_14; // @[TensorGemm.scala 346:19:@21410.4]
  assign mvc_io_wgt_data_bits_14_15 = io_wgt_rd_data_bits_14_15; // @[TensorGemm.scala 346:19:@21411.4]
  assign mvc_io_wgt_data_bits_15_0 = io_wgt_rd_data_bits_15_0; // @[TensorGemm.scala 346:19:@21412.4]
  assign mvc_io_wgt_data_bits_15_1 = io_wgt_rd_data_bits_15_1; // @[TensorGemm.scala 346:19:@21413.4]
  assign mvc_io_wgt_data_bits_15_2 = io_wgt_rd_data_bits_15_2; // @[TensorGemm.scala 346:19:@21414.4]
  assign mvc_io_wgt_data_bits_15_3 = io_wgt_rd_data_bits_15_3; // @[TensorGemm.scala 346:19:@21415.4]
  assign mvc_io_wgt_data_bits_15_4 = io_wgt_rd_data_bits_15_4; // @[TensorGemm.scala 346:19:@21416.4]
  assign mvc_io_wgt_data_bits_15_5 = io_wgt_rd_data_bits_15_5; // @[TensorGemm.scala 346:19:@21417.4]
  assign mvc_io_wgt_data_bits_15_6 = io_wgt_rd_data_bits_15_6; // @[TensorGemm.scala 346:19:@21418.4]
  assign mvc_io_wgt_data_bits_15_7 = io_wgt_rd_data_bits_15_7; // @[TensorGemm.scala 346:19:@21419.4]
  assign mvc_io_wgt_data_bits_15_8 = io_wgt_rd_data_bits_15_8; // @[TensorGemm.scala 346:19:@21420.4]
  assign mvc_io_wgt_data_bits_15_9 = io_wgt_rd_data_bits_15_9; // @[TensorGemm.scala 346:19:@21421.4]
  assign mvc_io_wgt_data_bits_15_10 = io_wgt_rd_data_bits_15_10; // @[TensorGemm.scala 346:19:@21422.4]
  assign mvc_io_wgt_data_bits_15_11 = io_wgt_rd_data_bits_15_11; // @[TensorGemm.scala 346:19:@21423.4]
  assign mvc_io_wgt_data_bits_15_12 = io_wgt_rd_data_bits_15_12; // @[TensorGemm.scala 346:19:@21424.4]
  assign mvc_io_wgt_data_bits_15_13 = io_wgt_rd_data_bits_15_13; // @[TensorGemm.scala 346:19:@21425.4]
  assign mvc_io_wgt_data_bits_15_14 = io_wgt_rd_data_bits_15_14; // @[TensorGemm.scala 346:19:@21426.4]
  assign mvc_io_wgt_data_bits_15_15 = io_wgt_rd_data_bits_15_15; // @[TensorGemm.scala 346:19:@21427.4]
  assign mvc_io_acc_i_data_valid = io_acc_rd_data_valid; // @[TensorGemm.scala 347:21:@21445.4]
  assign mvc_io_acc_i_data_bits_0_0 = io_acc_rd_data_bits_0_0; // @[TensorGemm.scala 347:21:@21429.4]
  assign mvc_io_acc_i_data_bits_0_1 = io_acc_rd_data_bits_0_1; // @[TensorGemm.scala 347:21:@21430.4]
  assign mvc_io_acc_i_data_bits_0_2 = io_acc_rd_data_bits_0_2; // @[TensorGemm.scala 347:21:@21431.4]
  assign mvc_io_acc_i_data_bits_0_3 = io_acc_rd_data_bits_0_3; // @[TensorGemm.scala 347:21:@21432.4]
  assign mvc_io_acc_i_data_bits_0_4 = io_acc_rd_data_bits_0_4; // @[TensorGemm.scala 347:21:@21433.4]
  assign mvc_io_acc_i_data_bits_0_5 = io_acc_rd_data_bits_0_5; // @[TensorGemm.scala 347:21:@21434.4]
  assign mvc_io_acc_i_data_bits_0_6 = io_acc_rd_data_bits_0_6; // @[TensorGemm.scala 347:21:@21435.4]
  assign mvc_io_acc_i_data_bits_0_7 = io_acc_rd_data_bits_0_7; // @[TensorGemm.scala 347:21:@21436.4]
  assign mvc_io_acc_i_data_bits_0_8 = io_acc_rd_data_bits_0_8; // @[TensorGemm.scala 347:21:@21437.4]
  assign mvc_io_acc_i_data_bits_0_9 = io_acc_rd_data_bits_0_9; // @[TensorGemm.scala 347:21:@21438.4]
  assign mvc_io_acc_i_data_bits_0_10 = io_acc_rd_data_bits_0_10; // @[TensorGemm.scala 347:21:@21439.4]
  assign mvc_io_acc_i_data_bits_0_11 = io_acc_rd_data_bits_0_11; // @[TensorGemm.scala 347:21:@21440.4]
  assign mvc_io_acc_i_data_bits_0_12 = io_acc_rd_data_bits_0_12; // @[TensorGemm.scala 347:21:@21441.4]
  assign mvc_io_acc_i_data_bits_0_13 = io_acc_rd_data_bits_0_13; // @[TensorGemm.scala 347:21:@21442.4]
  assign mvc_io_acc_i_data_bits_0_14 = io_acc_rd_data_bits_0_14; // @[TensorGemm.scala 347:21:@21443.4]
  assign mvc_io_acc_i_data_bits_0_15 = io_acc_rd_data_bits_0_15; // @[TensorGemm.scala 347:21:@21444.4]
  assign wrpipe_clock = clock; // @[:@20645.4]
  assign wrpipe_reset = reset; // @[:@20646.4]
  assign wrpipe_io_enq_valid = _T_7689 & _T_7830; // @[TensorGemm.scala 322:23:@20862.4]
  assign wrpipe_io_enq_bits = uop_acc; // @[TensorGemm.scala 323:22:@20863.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  uop_idx = _RAND_1[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  uop_acc = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  uop_inp = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  uop_wgt = _RAND_4[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  cnt_o = _RAND_5[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  acc_o = _RAND_6[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inp_o = _RAND_7[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wgt_o = _RAND_8[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  cnt_i = _RAND_9[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  acc_i = _RAND_10[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  inp_i = _RAND_11[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wgt_i = _RAND_12[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_7713) begin
        if (io_start) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_7714) begin
          state <= 3'h2;
        end else begin
          if (_T_7715) begin
            state <= 3'h3;
          end else begin
            if (_T_7716) begin
              state <= 3'h4;
            end else begin
              if (_T_7717) begin
                if (_T_7734) begin
                  if (_T_7736) begin
                    state <= 3'h5;
                  end else begin
                    state <= 3'h0;
                  end
                end else begin
                  state <= 3'h1;
                end
              end else begin
                if (_T_7737) begin
                  if (_T_7688) begin
                    state <= 3'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_7762) begin
      uop_idx <= {{1'd0}, dec_uop_begin};
    end else begin
      if (_T_7765) begin
        uop_idx <= _T_7768;
      end
    end
    if (_T_7822) begin
      uop_acc <= _T_7824;
    end
    if (_T_7822) begin
      uop_inp <= _T_7826;
    end
    if (_T_7822) begin
      uop_wgt <= _T_7828;
    end
    if (_T_7740) begin
      cnt_o <= 14'h0;
    end else begin
      if (_T_7786) begin
        cnt_o <= _T_7789;
      end
    end
    if (_T_7740) begin
      acc_o <= 14'h0;
    end else begin
      if (_T_7786) begin
        acc_o <= _T_7791;
      end
    end
    if (_T_7740) begin
      inp_o <= 14'h0;
    end else begin
      if (_T_7786) begin
        inp_o <= _T_7793;
      end
    end
    if (_T_7740) begin
      wgt_o <= 14'h0;
    end else begin
      if (_T_7786) begin
        wgt_o <= _T_7795;
      end
    end
    if (_T_7740) begin
      cnt_i <= 14'h0;
    end else begin
      if (_T_7803) begin
        cnt_i <= 14'h0;
      end else begin
        if (_T_7761) begin
          cnt_i <= _T_7814;
        end
      end
    end
    if (_T_7740) begin
      acc_i <= 14'h0;
    end else begin
      if (_T_7803) begin
        acc_i <= acc_o;
      end else begin
        if (_T_7761) begin
          acc_i <= _T_7816;
        end
      end
    end
    if (_T_7740) begin
      inp_i <= 14'h0;
    end else begin
      if (_T_7803) begin
        inp_i <= inp_o;
      end else begin
        if (_T_7761) begin
          inp_i <= _T_7818;
        end
      end
    end
    if (_T_7740) begin
      wgt_i <= 14'h0;
    end else begin
      if (_T_7803) begin
        wgt_i <= wgt_o;
      end else begin
        if (_T_7761) begin
          wgt_i <= _T_7820;
        end
      end
    end
    if (_T_7740) begin
      inflight <= 5'h0;
    end else begin
      if (_T_7743) begin
        if (!(_T_7745)) begin
          if (_T_7744) begin
            inflight <= _T_7749;
          end else begin
            if (mvc_io_acc_o_data_valid) begin
              inflight <= _T_7753;
            end
          end
        end
      end
    end
  end
endmodule
module Alu( // @[:@21490.2]
  input  [2:0]  io_opcode, // @[:@21493.4]
  input  [31:0] io_a, // @[:@21493.4]
  input  [31:0] io_b, // @[:@21493.4]
  output [31:0] io_y // @[:@21493.4]
);
  wire [31:0] ub; // @[TensorAlu.scala 37:17:@21495.4]
  wire [4:0] _T_13; // @[TensorAlu.scala 39:14:@21496.4]
  wire [4:0] _T_14; // @[TensorAlu.scala 39:11:@21497.4]
  wire [5:0] _T_16; // @[TensorAlu.scala 39:29:@21498.4]
  wire [4:0] m; // @[TensorAlu.scala 39:29:@21499.4]
  wire  _T_17; // @[TensorAlu.scala 42:26:@21501.4]
  wire [31:0] fop_0; // @[TensorAlu.scala 42:20:@21502.4]
  wire [31:0] fop_1; // @[TensorAlu.scala 42:50:@21504.4]
  wire [32:0] _T_19; // @[TensorAlu.scala 43:10:@21505.4]
  wire [31:0] _T_20; // @[TensorAlu.scala 43:10:@21506.4]
  wire [31:0] fop_2; // @[TensorAlu.scala 43:10:@21507.4]
  wire [31:0] fop_3; // @[TensorAlu.scala 43:23:@21508.4]
  wire [62:0] _GEN_0; // @[TensorAlu.scala 43:34:@21509.4]
  wire [62:0] fop_4; // @[TensorAlu.scala 43:34:@21509.4]
  wire  _T_21; // @[Mux.scala 46:19:@21510.4]
  wire [62:0] _T_22; // @[Mux.scala 46:16:@21511.4]
  wire  _T_23; // @[Mux.scala 46:19:@21512.4]
  wire [62:0] _T_24; // @[Mux.scala 46:16:@21513.4]
  wire  _T_25; // @[Mux.scala 46:19:@21514.4]
  wire [62:0] _T_26; // @[Mux.scala 46:16:@21515.4]
  wire  _T_27; // @[Mux.scala 46:19:@21516.4]
  wire [62:0] _T_28; // @[Mux.scala 46:16:@21517.4]
  wire  _T_29; // @[Mux.scala 46:19:@21518.4]
  wire [62:0] _T_30; // @[Mux.scala 46:16:@21519.4]
  wire [31:0] _GEN_1; // @[TensorAlu.scala 46:8:@21520.4]
  assign ub = $unsigned(io_b); // @[TensorAlu.scala 37:17:@21495.4]
  assign _T_13 = ub[4:0]; // @[TensorAlu.scala 39:14:@21496.4]
  assign _T_14 = ~ _T_13; // @[TensorAlu.scala 39:11:@21497.4]
  assign _T_16 = _T_14 + 5'h1; // @[TensorAlu.scala 39:29:@21498.4]
  assign m = _T_14 + 5'h1; // @[TensorAlu.scala 39:29:@21499.4]
  assign _T_17 = $signed(io_a) < $signed(io_b); // @[TensorAlu.scala 42:26:@21501.4]
  assign fop_0 = _T_17 ? $signed(io_a) : $signed(io_b); // @[TensorAlu.scala 42:20:@21502.4]
  assign fop_1 = _T_17 ? $signed(io_b) : $signed(io_a); // @[TensorAlu.scala 42:50:@21504.4]
  assign _T_19 = $signed(io_a) + $signed(io_b); // @[TensorAlu.scala 43:10:@21505.4]
  assign _T_20 = $signed(io_a) + $signed(io_b); // @[TensorAlu.scala 43:10:@21506.4]
  assign fop_2 = $signed(_T_20); // @[TensorAlu.scala 43:10:@21507.4]
  assign fop_3 = $signed(io_a) >>> _T_13; // @[TensorAlu.scala 43:23:@21508.4]
  assign _GEN_0 = {{31{io_a[31]}},io_a}; // @[TensorAlu.scala 43:34:@21509.4]
  assign fop_4 = $signed(_GEN_0) << m; // @[TensorAlu.scala 43:34:@21509.4]
  assign _T_21 = 3'h4 == io_opcode; // @[Mux.scala 46:19:@21510.4]
  assign _T_22 = _T_21 ? $signed(fop_4) : $signed({{31{io_a[31]}},io_a}); // @[Mux.scala 46:16:@21511.4]
  assign _T_23 = 3'h3 == io_opcode; // @[Mux.scala 46:19:@21512.4]
  assign _T_24 = _T_23 ? $signed({{31{fop_3[31]}},fop_3}) : $signed(_T_22); // @[Mux.scala 46:16:@21513.4]
  assign _T_25 = 3'h2 == io_opcode; // @[Mux.scala 46:19:@21514.4]
  assign _T_26 = _T_25 ? $signed({{31{fop_2[31]}},fop_2}) : $signed(_T_24); // @[Mux.scala 46:16:@21515.4]
  assign _T_27 = 3'h1 == io_opcode; // @[Mux.scala 46:19:@21516.4]
  assign _T_28 = _T_27 ? $signed({{31{fop_1[31]}},fop_1}) : $signed(_T_26); // @[Mux.scala 46:16:@21517.4]
  assign _T_29 = 3'h0 == io_opcode; // @[Mux.scala 46:19:@21518.4]
  assign _T_30 = _T_29 ? $signed({{31{fop_0[31]}},fop_0}) : $signed(_T_28); // @[Mux.scala 46:16:@21519.4]
  assign _GEN_1 = _T_30[31:0]; // @[TensorAlu.scala 46:8:@21520.4]
  assign io_y = $signed(_GEN_1); // @[TensorAlu.scala 46:8:@21520.4]
endmodule
module AluReg( // @[:@21522.2]
  input         clock, // @[:@21523.4]
  input  [2:0]  io_opcode, // @[:@21525.4]
  input         io_a_valid, // @[:@21525.4]
  input  [31:0] io_a_bits, // @[:@21525.4]
  input         io_b_valid, // @[:@21525.4]
  input  [31:0] io_b_bits, // @[:@21525.4]
  output        io_y_valid, // @[:@21525.4]
  output [31:0] io_y_bits // @[:@21525.4]
);
  wire [2:0] alu_io_opcode; // @[TensorAlu.scala 57:19:@21527.4]
  wire [31:0] alu_io_a; // @[TensorAlu.scala 57:19:@21527.4]
  wire [31:0] alu_io_b; // @[TensorAlu.scala 57:19:@21527.4]
  wire [31:0] alu_io_y; // @[TensorAlu.scala 57:19:@21527.4]
  reg [31:0] rA; // @[Reg.scala 11:16:@21530.4]
  reg [31:0] _RAND_0;
  reg [31:0] rB; // @[Reg.scala 11:16:@21534.4]
  reg [31:0] _RAND_1;
  reg  valid; // @[TensorAlu.scala 60:22:@21538.4]
  reg [31:0] _RAND_2;
  Alu alu ( // @[TensorAlu.scala 57:19:@21527.4]
    .io_opcode(alu_io_opcode),
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_y(alu_io_y)
  );
  assign io_y_valid = valid; // @[TensorAlu.scala 69:14:@21545.4]
  assign io_y_bits = $unsigned(alu_io_y); // @[TensorAlu.scala 70:13:@21547.4]
  assign alu_io_opcode = io_opcode; // @[TensorAlu.scala 62:17:@21540.4]
  assign alu_io_a = $signed(rA); // @[TensorAlu.scala 65:12:@21542.4]
  assign alu_io_b = $signed(rB); // @[TensorAlu.scala 66:12:@21544.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rA = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rB = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_a_valid) begin
      rA <= io_a_bits;
    end
    if (io_b_valid) begin
      rB <= io_b_bits;
    end
    valid <= io_b_valid;
  end
endmodule
module AluVector( // @[:@22434.2]
  input         clock, // @[:@22435.4]
  input  [2:0]  io_opcode, // @[:@22437.4]
  input         io_acc_a_data_valid, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_0, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_1, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_2, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_3, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_4, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_5, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_6, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_7, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_8, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_9, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_10, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_11, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_12, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_13, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_14, // @[:@22437.4]
  input  [31:0] io_acc_a_data_bits_0_15, // @[:@22437.4]
  input         io_acc_b_data_valid, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_0, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_1, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_2, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_3, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_4, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_5, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_6, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_7, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_8, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_9, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_10, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_11, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_12, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_13, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_14, // @[:@22437.4]
  input  [31:0] io_acc_b_data_bits_0_15, // @[:@22437.4]
  output        io_acc_y_data_valid, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_0, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_1, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_2, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_3, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_4, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_5, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_6, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_7, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_8, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_9, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_10, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_11, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_12, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_13, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_14, // @[:@22437.4]
  output [31:0] io_acc_y_data_bits_0_15, // @[:@22437.4]
  output        io_out_data_valid, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_0, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_1, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_2, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_3, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_4, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_5, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_6, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_7, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_8, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_9, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_10, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_11, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_12, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_13, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_14, // @[:@22437.4]
  output [7:0]  io_out_data_bits_0_15 // @[:@22437.4]
);
  wire  f_0_clock; // @[TensorAlu.scala 83:36:@22439.4]
  wire [2:0] f_0_io_opcode; // @[TensorAlu.scala 83:36:@22439.4]
  wire  f_0_io_a_valid; // @[TensorAlu.scala 83:36:@22439.4]
  wire [31:0] f_0_io_a_bits; // @[TensorAlu.scala 83:36:@22439.4]
  wire  f_0_io_b_valid; // @[TensorAlu.scala 83:36:@22439.4]
  wire [31:0] f_0_io_b_bits; // @[TensorAlu.scala 83:36:@22439.4]
  wire  f_0_io_y_valid; // @[TensorAlu.scala 83:36:@22439.4]
  wire [31:0] f_0_io_y_bits; // @[TensorAlu.scala 83:36:@22439.4]
  wire  f_1_clock; // @[TensorAlu.scala 83:36:@22442.4]
  wire [2:0] f_1_io_opcode; // @[TensorAlu.scala 83:36:@22442.4]
  wire  f_1_io_a_valid; // @[TensorAlu.scala 83:36:@22442.4]
  wire [31:0] f_1_io_a_bits; // @[TensorAlu.scala 83:36:@22442.4]
  wire  f_1_io_b_valid; // @[TensorAlu.scala 83:36:@22442.4]
  wire [31:0] f_1_io_b_bits; // @[TensorAlu.scala 83:36:@22442.4]
  wire  f_1_io_y_valid; // @[TensorAlu.scala 83:36:@22442.4]
  wire [31:0] f_1_io_y_bits; // @[TensorAlu.scala 83:36:@22442.4]
  wire  f_2_clock; // @[TensorAlu.scala 83:36:@22445.4]
  wire [2:0] f_2_io_opcode; // @[TensorAlu.scala 83:36:@22445.4]
  wire  f_2_io_a_valid; // @[TensorAlu.scala 83:36:@22445.4]
  wire [31:0] f_2_io_a_bits; // @[TensorAlu.scala 83:36:@22445.4]
  wire  f_2_io_b_valid; // @[TensorAlu.scala 83:36:@22445.4]
  wire [31:0] f_2_io_b_bits; // @[TensorAlu.scala 83:36:@22445.4]
  wire  f_2_io_y_valid; // @[TensorAlu.scala 83:36:@22445.4]
  wire [31:0] f_2_io_y_bits; // @[TensorAlu.scala 83:36:@22445.4]
  wire  f_3_clock; // @[TensorAlu.scala 83:36:@22448.4]
  wire [2:0] f_3_io_opcode; // @[TensorAlu.scala 83:36:@22448.4]
  wire  f_3_io_a_valid; // @[TensorAlu.scala 83:36:@22448.4]
  wire [31:0] f_3_io_a_bits; // @[TensorAlu.scala 83:36:@22448.4]
  wire  f_3_io_b_valid; // @[TensorAlu.scala 83:36:@22448.4]
  wire [31:0] f_3_io_b_bits; // @[TensorAlu.scala 83:36:@22448.4]
  wire  f_3_io_y_valid; // @[TensorAlu.scala 83:36:@22448.4]
  wire [31:0] f_3_io_y_bits; // @[TensorAlu.scala 83:36:@22448.4]
  wire  f_4_clock; // @[TensorAlu.scala 83:36:@22451.4]
  wire [2:0] f_4_io_opcode; // @[TensorAlu.scala 83:36:@22451.4]
  wire  f_4_io_a_valid; // @[TensorAlu.scala 83:36:@22451.4]
  wire [31:0] f_4_io_a_bits; // @[TensorAlu.scala 83:36:@22451.4]
  wire  f_4_io_b_valid; // @[TensorAlu.scala 83:36:@22451.4]
  wire [31:0] f_4_io_b_bits; // @[TensorAlu.scala 83:36:@22451.4]
  wire  f_4_io_y_valid; // @[TensorAlu.scala 83:36:@22451.4]
  wire [31:0] f_4_io_y_bits; // @[TensorAlu.scala 83:36:@22451.4]
  wire  f_5_clock; // @[TensorAlu.scala 83:36:@22454.4]
  wire [2:0] f_5_io_opcode; // @[TensorAlu.scala 83:36:@22454.4]
  wire  f_5_io_a_valid; // @[TensorAlu.scala 83:36:@22454.4]
  wire [31:0] f_5_io_a_bits; // @[TensorAlu.scala 83:36:@22454.4]
  wire  f_5_io_b_valid; // @[TensorAlu.scala 83:36:@22454.4]
  wire [31:0] f_5_io_b_bits; // @[TensorAlu.scala 83:36:@22454.4]
  wire  f_5_io_y_valid; // @[TensorAlu.scala 83:36:@22454.4]
  wire [31:0] f_5_io_y_bits; // @[TensorAlu.scala 83:36:@22454.4]
  wire  f_6_clock; // @[TensorAlu.scala 83:36:@22457.4]
  wire [2:0] f_6_io_opcode; // @[TensorAlu.scala 83:36:@22457.4]
  wire  f_6_io_a_valid; // @[TensorAlu.scala 83:36:@22457.4]
  wire [31:0] f_6_io_a_bits; // @[TensorAlu.scala 83:36:@22457.4]
  wire  f_6_io_b_valid; // @[TensorAlu.scala 83:36:@22457.4]
  wire [31:0] f_6_io_b_bits; // @[TensorAlu.scala 83:36:@22457.4]
  wire  f_6_io_y_valid; // @[TensorAlu.scala 83:36:@22457.4]
  wire [31:0] f_6_io_y_bits; // @[TensorAlu.scala 83:36:@22457.4]
  wire  f_7_clock; // @[TensorAlu.scala 83:36:@22460.4]
  wire [2:0] f_7_io_opcode; // @[TensorAlu.scala 83:36:@22460.4]
  wire  f_7_io_a_valid; // @[TensorAlu.scala 83:36:@22460.4]
  wire [31:0] f_7_io_a_bits; // @[TensorAlu.scala 83:36:@22460.4]
  wire  f_7_io_b_valid; // @[TensorAlu.scala 83:36:@22460.4]
  wire [31:0] f_7_io_b_bits; // @[TensorAlu.scala 83:36:@22460.4]
  wire  f_7_io_y_valid; // @[TensorAlu.scala 83:36:@22460.4]
  wire [31:0] f_7_io_y_bits; // @[TensorAlu.scala 83:36:@22460.4]
  wire  f_8_clock; // @[TensorAlu.scala 83:36:@22463.4]
  wire [2:0] f_8_io_opcode; // @[TensorAlu.scala 83:36:@22463.4]
  wire  f_8_io_a_valid; // @[TensorAlu.scala 83:36:@22463.4]
  wire [31:0] f_8_io_a_bits; // @[TensorAlu.scala 83:36:@22463.4]
  wire  f_8_io_b_valid; // @[TensorAlu.scala 83:36:@22463.4]
  wire [31:0] f_8_io_b_bits; // @[TensorAlu.scala 83:36:@22463.4]
  wire  f_8_io_y_valid; // @[TensorAlu.scala 83:36:@22463.4]
  wire [31:0] f_8_io_y_bits; // @[TensorAlu.scala 83:36:@22463.4]
  wire  f_9_clock; // @[TensorAlu.scala 83:36:@22466.4]
  wire [2:0] f_9_io_opcode; // @[TensorAlu.scala 83:36:@22466.4]
  wire  f_9_io_a_valid; // @[TensorAlu.scala 83:36:@22466.4]
  wire [31:0] f_9_io_a_bits; // @[TensorAlu.scala 83:36:@22466.4]
  wire  f_9_io_b_valid; // @[TensorAlu.scala 83:36:@22466.4]
  wire [31:0] f_9_io_b_bits; // @[TensorAlu.scala 83:36:@22466.4]
  wire  f_9_io_y_valid; // @[TensorAlu.scala 83:36:@22466.4]
  wire [31:0] f_9_io_y_bits; // @[TensorAlu.scala 83:36:@22466.4]
  wire  f_10_clock; // @[TensorAlu.scala 83:36:@22469.4]
  wire [2:0] f_10_io_opcode; // @[TensorAlu.scala 83:36:@22469.4]
  wire  f_10_io_a_valid; // @[TensorAlu.scala 83:36:@22469.4]
  wire [31:0] f_10_io_a_bits; // @[TensorAlu.scala 83:36:@22469.4]
  wire  f_10_io_b_valid; // @[TensorAlu.scala 83:36:@22469.4]
  wire [31:0] f_10_io_b_bits; // @[TensorAlu.scala 83:36:@22469.4]
  wire  f_10_io_y_valid; // @[TensorAlu.scala 83:36:@22469.4]
  wire [31:0] f_10_io_y_bits; // @[TensorAlu.scala 83:36:@22469.4]
  wire  f_11_clock; // @[TensorAlu.scala 83:36:@22472.4]
  wire [2:0] f_11_io_opcode; // @[TensorAlu.scala 83:36:@22472.4]
  wire  f_11_io_a_valid; // @[TensorAlu.scala 83:36:@22472.4]
  wire [31:0] f_11_io_a_bits; // @[TensorAlu.scala 83:36:@22472.4]
  wire  f_11_io_b_valid; // @[TensorAlu.scala 83:36:@22472.4]
  wire [31:0] f_11_io_b_bits; // @[TensorAlu.scala 83:36:@22472.4]
  wire  f_11_io_y_valid; // @[TensorAlu.scala 83:36:@22472.4]
  wire [31:0] f_11_io_y_bits; // @[TensorAlu.scala 83:36:@22472.4]
  wire  f_12_clock; // @[TensorAlu.scala 83:36:@22475.4]
  wire [2:0] f_12_io_opcode; // @[TensorAlu.scala 83:36:@22475.4]
  wire  f_12_io_a_valid; // @[TensorAlu.scala 83:36:@22475.4]
  wire [31:0] f_12_io_a_bits; // @[TensorAlu.scala 83:36:@22475.4]
  wire  f_12_io_b_valid; // @[TensorAlu.scala 83:36:@22475.4]
  wire [31:0] f_12_io_b_bits; // @[TensorAlu.scala 83:36:@22475.4]
  wire  f_12_io_y_valid; // @[TensorAlu.scala 83:36:@22475.4]
  wire [31:0] f_12_io_y_bits; // @[TensorAlu.scala 83:36:@22475.4]
  wire  f_13_clock; // @[TensorAlu.scala 83:36:@22478.4]
  wire [2:0] f_13_io_opcode; // @[TensorAlu.scala 83:36:@22478.4]
  wire  f_13_io_a_valid; // @[TensorAlu.scala 83:36:@22478.4]
  wire [31:0] f_13_io_a_bits; // @[TensorAlu.scala 83:36:@22478.4]
  wire  f_13_io_b_valid; // @[TensorAlu.scala 83:36:@22478.4]
  wire [31:0] f_13_io_b_bits; // @[TensorAlu.scala 83:36:@22478.4]
  wire  f_13_io_y_valid; // @[TensorAlu.scala 83:36:@22478.4]
  wire [31:0] f_13_io_y_bits; // @[TensorAlu.scala 83:36:@22478.4]
  wire  f_14_clock; // @[TensorAlu.scala 83:36:@22481.4]
  wire [2:0] f_14_io_opcode; // @[TensorAlu.scala 83:36:@22481.4]
  wire  f_14_io_a_valid; // @[TensorAlu.scala 83:36:@22481.4]
  wire [31:0] f_14_io_a_bits; // @[TensorAlu.scala 83:36:@22481.4]
  wire  f_14_io_b_valid; // @[TensorAlu.scala 83:36:@22481.4]
  wire [31:0] f_14_io_b_bits; // @[TensorAlu.scala 83:36:@22481.4]
  wire  f_14_io_y_valid; // @[TensorAlu.scala 83:36:@22481.4]
  wire [31:0] f_14_io_y_bits; // @[TensorAlu.scala 83:36:@22481.4]
  wire  f_15_clock; // @[TensorAlu.scala 83:36:@22484.4]
  wire [2:0] f_15_io_opcode; // @[TensorAlu.scala 83:36:@22484.4]
  wire  f_15_io_a_valid; // @[TensorAlu.scala 83:36:@22484.4]
  wire [31:0] f_15_io_a_bits; // @[TensorAlu.scala 83:36:@22484.4]
  wire  f_15_io_b_valid; // @[TensorAlu.scala 83:36:@22484.4]
  wire [31:0] f_15_io_b_bits; // @[TensorAlu.scala 83:36:@22484.4]
  wire  f_15_io_y_valid; // @[TensorAlu.scala 83:36:@22484.4]
  wire [31:0] f_15_io_y_bits; // @[TensorAlu.scala 83:36:@22484.4]
  wire  valid_1; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22501.4]
  wire  valid_0; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22493.4]
  wire  valid_3; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22517.4]
  wire  valid_2; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22509.4]
  wire  valid_5; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22533.4]
  wire  valid_4; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22525.4]
  wire  valid_7; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22549.4]
  wire  valid_6; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22541.4]
  wire [7:0] _T_1686; // @[TensorAlu.scala 95:32:@22622.4]
  wire  valid_9; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22565.4]
  wire  valid_8; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22557.4]
  wire  valid_11; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22581.4]
  wire  valid_10; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22573.4]
  wire  valid_13; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22597.4]
  wire  valid_12; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22589.4]
  wire  valid_15; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22613.4]
  wire  valid_14; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22605.4]
  wire [15:0] _T_1694; // @[TensorAlu.scala 95:32:@22630.4]
  wire [15:0] _T_1695; // @[TensorAlu.scala 95:39:@22631.4]
  AluReg f_0 ( // @[TensorAlu.scala 83:36:@22439.4]
    .clock(f_0_clock),
    .io_opcode(f_0_io_opcode),
    .io_a_valid(f_0_io_a_valid),
    .io_a_bits(f_0_io_a_bits),
    .io_b_valid(f_0_io_b_valid),
    .io_b_bits(f_0_io_b_bits),
    .io_y_valid(f_0_io_y_valid),
    .io_y_bits(f_0_io_y_bits)
  );
  AluReg f_1 ( // @[TensorAlu.scala 83:36:@22442.4]
    .clock(f_1_clock),
    .io_opcode(f_1_io_opcode),
    .io_a_valid(f_1_io_a_valid),
    .io_a_bits(f_1_io_a_bits),
    .io_b_valid(f_1_io_b_valid),
    .io_b_bits(f_1_io_b_bits),
    .io_y_valid(f_1_io_y_valid),
    .io_y_bits(f_1_io_y_bits)
  );
  AluReg f_2 ( // @[TensorAlu.scala 83:36:@22445.4]
    .clock(f_2_clock),
    .io_opcode(f_2_io_opcode),
    .io_a_valid(f_2_io_a_valid),
    .io_a_bits(f_2_io_a_bits),
    .io_b_valid(f_2_io_b_valid),
    .io_b_bits(f_2_io_b_bits),
    .io_y_valid(f_2_io_y_valid),
    .io_y_bits(f_2_io_y_bits)
  );
  AluReg f_3 ( // @[TensorAlu.scala 83:36:@22448.4]
    .clock(f_3_clock),
    .io_opcode(f_3_io_opcode),
    .io_a_valid(f_3_io_a_valid),
    .io_a_bits(f_3_io_a_bits),
    .io_b_valid(f_3_io_b_valid),
    .io_b_bits(f_3_io_b_bits),
    .io_y_valid(f_3_io_y_valid),
    .io_y_bits(f_3_io_y_bits)
  );
  AluReg f_4 ( // @[TensorAlu.scala 83:36:@22451.4]
    .clock(f_4_clock),
    .io_opcode(f_4_io_opcode),
    .io_a_valid(f_4_io_a_valid),
    .io_a_bits(f_4_io_a_bits),
    .io_b_valid(f_4_io_b_valid),
    .io_b_bits(f_4_io_b_bits),
    .io_y_valid(f_4_io_y_valid),
    .io_y_bits(f_4_io_y_bits)
  );
  AluReg f_5 ( // @[TensorAlu.scala 83:36:@22454.4]
    .clock(f_5_clock),
    .io_opcode(f_5_io_opcode),
    .io_a_valid(f_5_io_a_valid),
    .io_a_bits(f_5_io_a_bits),
    .io_b_valid(f_5_io_b_valid),
    .io_b_bits(f_5_io_b_bits),
    .io_y_valid(f_5_io_y_valid),
    .io_y_bits(f_5_io_y_bits)
  );
  AluReg f_6 ( // @[TensorAlu.scala 83:36:@22457.4]
    .clock(f_6_clock),
    .io_opcode(f_6_io_opcode),
    .io_a_valid(f_6_io_a_valid),
    .io_a_bits(f_6_io_a_bits),
    .io_b_valid(f_6_io_b_valid),
    .io_b_bits(f_6_io_b_bits),
    .io_y_valid(f_6_io_y_valid),
    .io_y_bits(f_6_io_y_bits)
  );
  AluReg f_7 ( // @[TensorAlu.scala 83:36:@22460.4]
    .clock(f_7_clock),
    .io_opcode(f_7_io_opcode),
    .io_a_valid(f_7_io_a_valid),
    .io_a_bits(f_7_io_a_bits),
    .io_b_valid(f_7_io_b_valid),
    .io_b_bits(f_7_io_b_bits),
    .io_y_valid(f_7_io_y_valid),
    .io_y_bits(f_7_io_y_bits)
  );
  AluReg f_8 ( // @[TensorAlu.scala 83:36:@22463.4]
    .clock(f_8_clock),
    .io_opcode(f_8_io_opcode),
    .io_a_valid(f_8_io_a_valid),
    .io_a_bits(f_8_io_a_bits),
    .io_b_valid(f_8_io_b_valid),
    .io_b_bits(f_8_io_b_bits),
    .io_y_valid(f_8_io_y_valid),
    .io_y_bits(f_8_io_y_bits)
  );
  AluReg f_9 ( // @[TensorAlu.scala 83:36:@22466.4]
    .clock(f_9_clock),
    .io_opcode(f_9_io_opcode),
    .io_a_valid(f_9_io_a_valid),
    .io_a_bits(f_9_io_a_bits),
    .io_b_valid(f_9_io_b_valid),
    .io_b_bits(f_9_io_b_bits),
    .io_y_valid(f_9_io_y_valid),
    .io_y_bits(f_9_io_y_bits)
  );
  AluReg f_10 ( // @[TensorAlu.scala 83:36:@22469.4]
    .clock(f_10_clock),
    .io_opcode(f_10_io_opcode),
    .io_a_valid(f_10_io_a_valid),
    .io_a_bits(f_10_io_a_bits),
    .io_b_valid(f_10_io_b_valid),
    .io_b_bits(f_10_io_b_bits),
    .io_y_valid(f_10_io_y_valid),
    .io_y_bits(f_10_io_y_bits)
  );
  AluReg f_11 ( // @[TensorAlu.scala 83:36:@22472.4]
    .clock(f_11_clock),
    .io_opcode(f_11_io_opcode),
    .io_a_valid(f_11_io_a_valid),
    .io_a_bits(f_11_io_a_bits),
    .io_b_valid(f_11_io_b_valid),
    .io_b_bits(f_11_io_b_bits),
    .io_y_valid(f_11_io_y_valid),
    .io_y_bits(f_11_io_y_bits)
  );
  AluReg f_12 ( // @[TensorAlu.scala 83:36:@22475.4]
    .clock(f_12_clock),
    .io_opcode(f_12_io_opcode),
    .io_a_valid(f_12_io_a_valid),
    .io_a_bits(f_12_io_a_bits),
    .io_b_valid(f_12_io_b_valid),
    .io_b_bits(f_12_io_b_bits),
    .io_y_valid(f_12_io_y_valid),
    .io_y_bits(f_12_io_y_bits)
  );
  AluReg f_13 ( // @[TensorAlu.scala 83:36:@22478.4]
    .clock(f_13_clock),
    .io_opcode(f_13_io_opcode),
    .io_a_valid(f_13_io_a_valid),
    .io_a_bits(f_13_io_a_bits),
    .io_b_valid(f_13_io_b_valid),
    .io_b_bits(f_13_io_b_bits),
    .io_y_valid(f_13_io_y_valid),
    .io_y_bits(f_13_io_y_bits)
  );
  AluReg f_14 ( // @[TensorAlu.scala 83:36:@22481.4]
    .clock(f_14_clock),
    .io_opcode(f_14_io_opcode),
    .io_a_valid(f_14_io_a_valid),
    .io_a_bits(f_14_io_a_bits),
    .io_b_valid(f_14_io_b_valid),
    .io_b_bits(f_14_io_b_bits),
    .io_y_valid(f_14_io_y_valid),
    .io_y_bits(f_14_io_y_bits)
  );
  AluReg f_15 ( // @[TensorAlu.scala 83:36:@22484.4]
    .clock(f_15_clock),
    .io_opcode(f_15_io_opcode),
    .io_a_valid(f_15_io_a_valid),
    .io_a_bits(f_15_io_a_bits),
    .io_b_valid(f_15_io_b_valid),
    .io_b_bits(f_15_io_b_bits),
    .io_y_valid(f_15_io_y_valid),
    .io_y_bits(f_15_io_y_bits)
  );
  assign valid_1 = f_1_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22501.4]
  assign valid_0 = f_0_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22493.4]
  assign valid_3 = f_3_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22517.4]
  assign valid_2 = f_2_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22509.4]
  assign valid_5 = f_5_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22533.4]
  assign valid_4 = f_4_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22525.4]
  assign valid_7 = f_7_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22549.4]
  assign valid_6 = f_6_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22541.4]
  assign _T_1686 = {valid_7,valid_6,valid_5,valid_4,valid_3,valid_2,valid_1,valid_0}; // @[TensorAlu.scala 95:32:@22622.4]
  assign valid_9 = f_9_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22565.4]
  assign valid_8 = f_8_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22557.4]
  assign valid_11 = f_11_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22581.4]
  assign valid_10 = f_10_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22573.4]
  assign valid_13 = f_13_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22597.4]
  assign valid_12 = f_12_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22589.4]
  assign valid_15 = f_15_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22613.4]
  assign valid_14 = f_14_io_y_valid; // @[TensorAlu.scala 84:19:@22487.4 TensorAlu.scala 91:14:@22605.4]
  assign _T_1694 = {valid_15,valid_14,valid_13,valid_12,valid_11,valid_10,valid_9,valid_8,_T_1686}; // @[TensorAlu.scala 95:32:@22630.4]
  assign _T_1695 = ~ _T_1694; // @[TensorAlu.scala 95:39:@22631.4]
  assign io_acc_y_data_valid = _T_1695 == 16'h0; // @[TensorAlu.scala 95:23:@22633.4]
  assign io_acc_y_data_bits_0_0 = f_0_io_y_bits; // @[TensorAlu.scala 92:30:@22494.4]
  assign io_acc_y_data_bits_0_1 = f_1_io_y_bits; // @[TensorAlu.scala 92:30:@22502.4]
  assign io_acc_y_data_bits_0_2 = f_2_io_y_bits; // @[TensorAlu.scala 92:30:@22510.4]
  assign io_acc_y_data_bits_0_3 = f_3_io_y_bits; // @[TensorAlu.scala 92:30:@22518.4]
  assign io_acc_y_data_bits_0_4 = f_4_io_y_bits; // @[TensorAlu.scala 92:30:@22526.4]
  assign io_acc_y_data_bits_0_5 = f_5_io_y_bits; // @[TensorAlu.scala 92:30:@22534.4]
  assign io_acc_y_data_bits_0_6 = f_6_io_y_bits; // @[TensorAlu.scala 92:30:@22542.4]
  assign io_acc_y_data_bits_0_7 = f_7_io_y_bits; // @[TensorAlu.scala 92:30:@22550.4]
  assign io_acc_y_data_bits_0_8 = f_8_io_y_bits; // @[TensorAlu.scala 92:30:@22558.4]
  assign io_acc_y_data_bits_0_9 = f_9_io_y_bits; // @[TensorAlu.scala 92:30:@22566.4]
  assign io_acc_y_data_bits_0_10 = f_10_io_y_bits; // @[TensorAlu.scala 92:30:@22574.4]
  assign io_acc_y_data_bits_0_11 = f_11_io_y_bits; // @[TensorAlu.scala 92:30:@22582.4]
  assign io_acc_y_data_bits_0_12 = f_12_io_y_bits; // @[TensorAlu.scala 92:30:@22590.4]
  assign io_acc_y_data_bits_0_13 = f_13_io_y_bits; // @[TensorAlu.scala 92:30:@22598.4]
  assign io_acc_y_data_bits_0_14 = f_14_io_y_bits; // @[TensorAlu.scala 92:30:@22606.4]
  assign io_acc_y_data_bits_0_15 = f_15_io_y_bits; // @[TensorAlu.scala 92:30:@22614.4]
  assign io_out_data_valid = _T_1695 == 16'h0; // @[TensorAlu.scala 96:21:@22651.4]
  assign io_out_data_bits_0_0 = f_0_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22495.4]
  assign io_out_data_bits_0_1 = f_1_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22503.4]
  assign io_out_data_bits_0_2 = f_2_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22511.4]
  assign io_out_data_bits_0_3 = f_3_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22519.4]
  assign io_out_data_bits_0_4 = f_4_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22527.4]
  assign io_out_data_bits_0_5 = f_5_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22535.4]
  assign io_out_data_bits_0_6 = f_6_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22543.4]
  assign io_out_data_bits_0_7 = f_7_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22551.4]
  assign io_out_data_bits_0_8 = f_8_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22559.4]
  assign io_out_data_bits_0_9 = f_9_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22567.4]
  assign io_out_data_bits_0_10 = f_10_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22575.4]
  assign io_out_data_bits_0_11 = f_11_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22583.4]
  assign io_out_data_bits_0_12 = f_12_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22591.4]
  assign io_out_data_bits_0_13 = f_13_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22599.4]
  assign io_out_data_bits_0_14 = f_14_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22607.4]
  assign io_out_data_bits_0_15 = f_15_io_y_bits[7:0]; // @[TensorAlu.scala 93:28:@22615.4]
  assign f_0_clock = clock; // @[:@22440.4]
  assign f_0_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22488.4]
  assign f_0_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22489.4]
  assign f_0_io_a_bits = io_acc_a_data_bits_0_0; // @[TensorAlu.scala 88:20:@22490.4]
  assign f_0_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22491.4]
  assign f_0_io_b_bits = io_acc_b_data_bits_0_0; // @[TensorAlu.scala 90:20:@22492.4]
  assign f_1_clock = clock; // @[:@22443.4]
  assign f_1_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22496.4]
  assign f_1_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22497.4]
  assign f_1_io_a_bits = io_acc_a_data_bits_0_1; // @[TensorAlu.scala 88:20:@22498.4]
  assign f_1_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22499.4]
  assign f_1_io_b_bits = io_acc_b_data_bits_0_1; // @[TensorAlu.scala 90:20:@22500.4]
  assign f_2_clock = clock; // @[:@22446.4]
  assign f_2_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22504.4]
  assign f_2_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22505.4]
  assign f_2_io_a_bits = io_acc_a_data_bits_0_2; // @[TensorAlu.scala 88:20:@22506.4]
  assign f_2_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22507.4]
  assign f_2_io_b_bits = io_acc_b_data_bits_0_2; // @[TensorAlu.scala 90:20:@22508.4]
  assign f_3_clock = clock; // @[:@22449.4]
  assign f_3_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22512.4]
  assign f_3_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22513.4]
  assign f_3_io_a_bits = io_acc_a_data_bits_0_3; // @[TensorAlu.scala 88:20:@22514.4]
  assign f_3_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22515.4]
  assign f_3_io_b_bits = io_acc_b_data_bits_0_3; // @[TensorAlu.scala 90:20:@22516.4]
  assign f_4_clock = clock; // @[:@22452.4]
  assign f_4_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22520.4]
  assign f_4_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22521.4]
  assign f_4_io_a_bits = io_acc_a_data_bits_0_4; // @[TensorAlu.scala 88:20:@22522.4]
  assign f_4_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22523.4]
  assign f_4_io_b_bits = io_acc_b_data_bits_0_4; // @[TensorAlu.scala 90:20:@22524.4]
  assign f_5_clock = clock; // @[:@22455.4]
  assign f_5_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22528.4]
  assign f_5_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22529.4]
  assign f_5_io_a_bits = io_acc_a_data_bits_0_5; // @[TensorAlu.scala 88:20:@22530.4]
  assign f_5_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22531.4]
  assign f_5_io_b_bits = io_acc_b_data_bits_0_5; // @[TensorAlu.scala 90:20:@22532.4]
  assign f_6_clock = clock; // @[:@22458.4]
  assign f_6_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22536.4]
  assign f_6_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22537.4]
  assign f_6_io_a_bits = io_acc_a_data_bits_0_6; // @[TensorAlu.scala 88:20:@22538.4]
  assign f_6_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22539.4]
  assign f_6_io_b_bits = io_acc_b_data_bits_0_6; // @[TensorAlu.scala 90:20:@22540.4]
  assign f_7_clock = clock; // @[:@22461.4]
  assign f_7_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22544.4]
  assign f_7_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22545.4]
  assign f_7_io_a_bits = io_acc_a_data_bits_0_7; // @[TensorAlu.scala 88:20:@22546.4]
  assign f_7_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22547.4]
  assign f_7_io_b_bits = io_acc_b_data_bits_0_7; // @[TensorAlu.scala 90:20:@22548.4]
  assign f_8_clock = clock; // @[:@22464.4]
  assign f_8_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22552.4]
  assign f_8_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22553.4]
  assign f_8_io_a_bits = io_acc_a_data_bits_0_8; // @[TensorAlu.scala 88:20:@22554.4]
  assign f_8_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22555.4]
  assign f_8_io_b_bits = io_acc_b_data_bits_0_8; // @[TensorAlu.scala 90:20:@22556.4]
  assign f_9_clock = clock; // @[:@22467.4]
  assign f_9_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22560.4]
  assign f_9_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22561.4]
  assign f_9_io_a_bits = io_acc_a_data_bits_0_9; // @[TensorAlu.scala 88:20:@22562.4]
  assign f_9_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22563.4]
  assign f_9_io_b_bits = io_acc_b_data_bits_0_9; // @[TensorAlu.scala 90:20:@22564.4]
  assign f_10_clock = clock; // @[:@22470.4]
  assign f_10_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22568.4]
  assign f_10_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22569.4]
  assign f_10_io_a_bits = io_acc_a_data_bits_0_10; // @[TensorAlu.scala 88:20:@22570.4]
  assign f_10_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22571.4]
  assign f_10_io_b_bits = io_acc_b_data_bits_0_10; // @[TensorAlu.scala 90:20:@22572.4]
  assign f_11_clock = clock; // @[:@22473.4]
  assign f_11_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22576.4]
  assign f_11_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22577.4]
  assign f_11_io_a_bits = io_acc_a_data_bits_0_11; // @[TensorAlu.scala 88:20:@22578.4]
  assign f_11_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22579.4]
  assign f_11_io_b_bits = io_acc_b_data_bits_0_11; // @[TensorAlu.scala 90:20:@22580.4]
  assign f_12_clock = clock; // @[:@22476.4]
  assign f_12_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22584.4]
  assign f_12_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22585.4]
  assign f_12_io_a_bits = io_acc_a_data_bits_0_12; // @[TensorAlu.scala 88:20:@22586.4]
  assign f_12_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22587.4]
  assign f_12_io_b_bits = io_acc_b_data_bits_0_12; // @[TensorAlu.scala 90:20:@22588.4]
  assign f_13_clock = clock; // @[:@22479.4]
  assign f_13_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22592.4]
  assign f_13_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22593.4]
  assign f_13_io_a_bits = io_acc_a_data_bits_0_13; // @[TensorAlu.scala 88:20:@22594.4]
  assign f_13_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22595.4]
  assign f_13_io_b_bits = io_acc_b_data_bits_0_13; // @[TensorAlu.scala 90:20:@22596.4]
  assign f_14_clock = clock; // @[:@22482.4]
  assign f_14_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22600.4]
  assign f_14_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22601.4]
  assign f_14_io_a_bits = io_acc_a_data_bits_0_14; // @[TensorAlu.scala 88:20:@22602.4]
  assign f_14_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22603.4]
  assign f_14_io_b_bits = io_acc_b_data_bits_0_14; // @[TensorAlu.scala 90:20:@22604.4]
  assign f_15_clock = clock; // @[:@22485.4]
  assign f_15_io_opcode = io_opcode; // @[TensorAlu.scala 86:20:@22608.4]
  assign f_15_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 87:21:@22609.4]
  assign f_15_io_a_bits = io_acc_a_data_bits_0_15; // @[TensorAlu.scala 88:20:@22610.4]
  assign f_15_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 89:21:@22611.4]
  assign f_15_io_b_bits = io_acc_b_data_bits_0_15; // @[TensorAlu.scala 90:20:@22612.4]
endmodule
module TensorAlu( // @[:@22653.2]
  input          clock, // @[:@22654.4]
  input          reset, // @[:@22655.4]
  input          io_start, // @[:@22656.4]
  output         io_done, // @[:@22656.4]
  input  [127:0] io_inst, // @[:@22656.4]
  output         io_uop_idx_valid, // @[:@22656.4]
  output [10:0]  io_uop_idx_bits, // @[:@22656.4]
  input          io_uop_data_valid, // @[:@22656.4]
  input  [10:0]  io_uop_data_bits_u1, // @[:@22656.4]
  input  [10:0]  io_uop_data_bits_u0, // @[:@22656.4]
  output         io_acc_rd_idx_valid, // @[:@22656.4]
  output [10:0]  io_acc_rd_idx_bits, // @[:@22656.4]
  input          io_acc_rd_data_valid, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_0, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_1, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_2, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_3, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_4, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_5, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_6, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_7, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_8, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_9, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_10, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_11, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_12, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_13, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_14, // @[:@22656.4]
  input  [31:0]  io_acc_rd_data_bits_0_15, // @[:@22656.4]
  output         io_acc_wr_valid, // @[:@22656.4]
  output [10:0]  io_acc_wr_bits_idx, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_0, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_1, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_2, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_3, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_4, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_5, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_6, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_7, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_8, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_9, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_10, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_11, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_12, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_13, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_14, // @[:@22656.4]
  output [31:0]  io_acc_wr_bits_data_0_15, // @[:@22656.4]
  output         io_out_wr_valid, // @[:@22656.4]
  output [10:0]  io_out_wr_bits_idx, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_0, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_1, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_2, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_3, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_4, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_5, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_6, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_7, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_8, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_9, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_10, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_11, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_12, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_13, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_14, // @[:@22656.4]
  output [7:0]   io_out_wr_bits_data_0_15 // @[:@22656.4]
);
  wire  alu_clock; // @[TensorAlu.scala 119:19:@22659.4]
  wire [2:0] alu_io_opcode; // @[TensorAlu.scala 119:19:@22659.4]
  wire  alu_io_acc_a_data_valid; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_0; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_1; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_2; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_3; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_4; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_5; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_6; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_7; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_8; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_9; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_10; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_11; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_12; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_13; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_14; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_a_data_bits_0_15; // @[TensorAlu.scala 119:19:@22659.4]
  wire  alu_io_acc_b_data_valid; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_0; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_1; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_2; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_3; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_4; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_5; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_6; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_7; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_8; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_9; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_10; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_11; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_12; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_13; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_14; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_b_data_bits_0_15; // @[TensorAlu.scala 119:19:@22659.4]
  wire  alu_io_acc_y_data_valid; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_0; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_1; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_2; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_3; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_4; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_5; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_6; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_7; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_8; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_9; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_10; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_11; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_12; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_13; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_14; // @[TensorAlu.scala 119:19:@22659.4]
  wire [31:0] alu_io_acc_y_data_bits_0_15; // @[TensorAlu.scala 119:19:@22659.4]
  wire  alu_io_out_data_valid; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_0; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_1; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_2; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_3; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_4; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_5; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_6; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_7; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_8; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_9; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_10; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_11; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_12; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_13; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_14; // @[TensorAlu.scala 119:19:@22659.4]
  wire [7:0] alu_io_out_data_bits_0_15; // @[TensorAlu.scala 119:19:@22659.4]
  reg [2:0] state; // @[TensorAlu.scala 118:22:@22658.4]
  reg [31:0] _RAND_0;
  wire [12:0] dec_uop_begin; // @[TensorAlu.scala 120:29:@22677.4]
  wire [13:0] dec_uop_end; // @[TensorAlu.scala 120:29:@22679.4]
  wire [13:0] dec_lp_0; // @[TensorAlu.scala 120:29:@22681.4]
  wire [13:0] dec_lp_1; // @[TensorAlu.scala 120:29:@22683.4]
  wire [10:0] dec_dst_0; // @[TensorAlu.scala 120:29:@22687.4]
  wire [10:0] dec_dst_1; // @[TensorAlu.scala 120:29:@22689.4]
  wire [10:0] dec_src_0; // @[TensorAlu.scala 120:29:@22691.4]
  wire [10:0] dec_src_1; // @[TensorAlu.scala 120:29:@22693.4]
  wire [1:0] dec_alu_op; // @[TensorAlu.scala 120:29:@22695.4]
  wire  dec_alu_use_imm; // @[TensorAlu.scala 120:29:@22697.4]
  wire [15:0] dec_alu_imm; // @[TensorAlu.scala 120:29:@22699.4]
  reg [13:0] uop_idx; // @[TensorAlu.scala 121:20:@22703.4]
  reg [31:0] _RAND_1;
  reg [13:0] uop_dst; // @[TensorAlu.scala 123:20:@22704.4]
  reg [31:0] _RAND_2;
  reg [13:0] uop_src; // @[TensorAlu.scala 124:20:@22705.4]
  reg [31:0] _RAND_3;
  reg [13:0] cnt_o; // @[TensorAlu.scala 125:18:@22706.4]
  reg [31:0] _RAND_4;
  reg [13:0] dst_o; // @[TensorAlu.scala 126:18:@22707.4]
  reg [31:0] _RAND_5;
  reg [13:0] src_o; // @[TensorAlu.scala 127:18:@22708.4]
  reg [31:0] _RAND_6;
  reg [13:0] cnt_i; // @[TensorAlu.scala 128:18:@22709.4]
  reg [31:0] _RAND_7;
  reg [13:0] dst_i; // @[TensorAlu.scala 129:18:@22710.4]
  reg [31:0] _RAND_8;
  reg [13:0] src_i; // @[TensorAlu.scala 130:18:@22711.4]
  reg [31:0] _RAND_9;
  wire  _T_1440; // @[TensorAlu.scala 132:11:@22712.4]
  wire  _T_1441; // @[TensorAlu.scala 132:20:@22713.4]
  wire [14:0] _T_1443; // @[TensorAlu.scala 134:27:@22714.4]
  wire [14:0] _T_1444; // @[TensorAlu.scala 134:27:@22715.4]
  wire [13:0] _T_1445; // @[TensorAlu.scala 134:27:@22716.4]
  wire  _T_1446; // @[TensorAlu.scala 134:14:@22717.4]
  wire  _T_1447; // @[TensorAlu.scala 133:29:@22718.4]
  wire [14:0] _T_1449; // @[TensorAlu.scala 135:27:@22719.4]
  wire [14:0] _T_1450; // @[TensorAlu.scala 135:27:@22720.4]
  wire [13:0] _T_1451; // @[TensorAlu.scala 135:27:@22721.4]
  wire  _T_1452; // @[TensorAlu.scala 135:14:@22722.4]
  wire  _T_1453; // @[TensorAlu.scala 134:34:@22723.4]
  wire [14:0] _T_1455; // @[TensorAlu.scala 136:28:@22724.4]
  wire [14:0] _T_1456; // @[TensorAlu.scala 136:28:@22725.4]
  wire [13:0] _T_1457; // @[TensorAlu.scala 136:28:@22726.4]
  wire  _T_1458; // @[TensorAlu.scala 136:16:@22727.4]
  wire  _T_1459; // @[Conditional.scala 37:30:@22729.4]
  wire [2:0] _GEN_0; // @[TensorAlu.scala 140:22:@22731.6]
  wire  _T_1460; // @[Conditional.scala 37:30:@22736.6]
  wire  _T_1461; // @[Conditional.scala 37:30:@22741.8]
  wire  _T_1462; // @[Conditional.scala 37:30:@22746.10]
  wire  _T_1463; // @[Conditional.scala 37:30:@22751.12]
  wire  _T_1464; // @[Conditional.scala 37:30:@22756.14]
  wire  _T_1475; // @[TensorAlu.scala 159:38:@22767.18]
  wire  _T_1481; // @[TensorAlu.scala 160:40:@22772.18]
  wire [2:0] _GEN_1; // @[TensorAlu.scala 161:42:@22773.18]
  wire [2:0] _GEN_2; // @[TensorAlu.scala 157:35:@22758.16]
  wire [2:0] _GEN_3; // @[Conditional.scala 39:67:@22757.14]
  wire [2:0] _GEN_4; // @[Conditional.scala 39:67:@22752.12]
  wire [2:0] _GEN_5; // @[Conditional.scala 39:67:@22747.10]
  wire [2:0] _GEN_6; // @[Conditional.scala 39:67:@22742.8]
  wire [2:0] _GEN_7; // @[Conditional.scala 39:67:@22737.6]
  wire [2:0] _GEN_8; // @[Conditional.scala 40:58:@22730.4]
  wire  _T_1482; // @[TensorAlu.scala 171:11:@22781.4]
  wire  _T_1490; // @[TensorAlu.scala 173:31:@22788.4]
  wire  _T_1491; // @[TensorAlu.scala 171:21:@22789.4]
  wire [14:0] _T_1495; // @[TensorAlu.scala 177:24:@22797.8]
  wire [13:0] _T_1496; // @[TensorAlu.scala 177:24:@22798.8]
  wire [13:0] _GEN_9; // @[TensorAlu.scala 176:55:@22796.6]
  wire  _T_1514; // @[TensorAlu.scala 187:33:@22819.6]
  wire [14:0] _T_1516; // @[TensorAlu.scala 189:20:@22821.8]
  wire [13:0] _T_1517; // @[TensorAlu.scala 189:20:@22822.8]
  wire [13:0] _GEN_28; // @[TensorAlu.scala 190:20:@22824.8]
  wire [14:0] _T_1518; // @[TensorAlu.scala 190:20:@22824.8]
  wire [13:0] _T_1519; // @[TensorAlu.scala 190:20:@22825.8]
  wire [13:0] _GEN_29; // @[TensorAlu.scala 191:20:@22827.8]
  wire [14:0] _T_1520; // @[TensorAlu.scala 191:20:@22827.8]
  wire [13:0] _T_1521; // @[TensorAlu.scala 191:20:@22828.8]
  wire [13:0] _GEN_11; // @[TensorAlu.scala 188:33:@22820.6]
  wire [13:0] _GEN_12; // @[TensorAlu.scala 188:33:@22820.6]
  wire [13:0] _GEN_13; // @[TensorAlu.scala 188:33:@22820.6]
  wire  _T_1526; // @[TensorAlu.scala 198:20:@22838.6]
  wire  _T_1527; // @[TensorAlu.scala 198:42:@22839.6]
  wire  _T_1528; // @[TensorAlu.scala 198:33:@22840.6]
  wire [14:0] _T_1539; // @[TensorAlu.scala 203:20:@22855.10]
  wire [13:0] _T_1540; // @[TensorAlu.scala 203:20:@22856.10]
  wire [13:0] _GEN_30; // @[TensorAlu.scala 204:20:@22858.10]
  wire [14:0] _T_1541; // @[TensorAlu.scala 204:20:@22858.10]
  wire [13:0] _T_1542; // @[TensorAlu.scala 204:20:@22859.10]
  wire [13:0] _GEN_31; // @[TensorAlu.scala 205:20:@22861.10]
  wire [14:0] _T_1543; // @[TensorAlu.scala 205:20:@22861.10]
  wire [13:0] _T_1544; // @[TensorAlu.scala 205:20:@22862.10]
  wire [13:0] _GEN_17; // @[TensorAlu.scala 202:84:@22854.8]
  wire [13:0] _GEN_18; // @[TensorAlu.scala 202:84:@22854.8]
  wire [13:0] _GEN_19; // @[TensorAlu.scala 202:84:@22854.8]
  wire [13:0] _GEN_20; // @[TensorAlu.scala 198:56:@22841.6]
  wire [13:0] _GEN_21; // @[TensorAlu.scala 198:56:@22841.6]
  wire [13:0] _GEN_22; // @[TensorAlu.scala 198:56:@22841.6]
  wire  _T_1545; // @[TensorAlu.scala 208:14:@22865.4]
  wire  _T_1546; // @[TensorAlu.scala 208:30:@22866.4]
  wire [13:0] _GEN_32; // @[TensorAlu.scala 209:36:@22868.6]
  wire [14:0] _T_1547; // @[TensorAlu.scala 209:36:@22868.6]
  wire [13:0] _T_1548; // @[TensorAlu.scala 209:36:@22869.6]
  wire [13:0] _GEN_33; // @[TensorAlu.scala 210:36:@22871.6]
  wire [14:0] _T_1549; // @[TensorAlu.scala 210:36:@22871.6]
  wire [13:0] _T_1550; // @[TensorAlu.scala 210:36:@22872.6]
  wire  _T_1552; // @[TensorAlu.scala 218:32:@22878.4]
  wire  _T_1553; // @[TensorAlu.scala 218:58:@22879.4]
  wire  _T_1554; // @[TensorAlu.scala 218:77:@22880.4]
  wire  _T_1555; // @[TensorAlu.scala 218:75:@22881.4]
  wire [13:0] _T_1558; // @[TensorAlu.scala 219:28:@22885.4]
  wire  _T_1863; // @[TensorAlu.scala 226:27:@22890.4]
  wire [31:0] _T_1866; // @[Cat.scala 30:58:@22892.4]
  wire [31:0] tensorImm_data_bits_0_0; // @[TensorAlu.scala 226:15:@22893.4]
  wire [2:0] _GEN_34; // @[TensorAlu.scala 232:26:@22970.4]
  wire  isSHR; // @[TensorAlu.scala 232:26:@22970.4]
  wire  neg_shift; // @[TensorAlu.scala 233:25:@22972.4]
  wire [1:0] _T_1945; // @[TensorAlu.scala 234:40:@22973.4]
  wire  _T_1949; // @[TensorAlu.scala 240:26:@22996.4]
  AluVector alu ( // @[TensorAlu.scala 119:19:@22659.4]
    .clock(alu_clock),
    .io_opcode(alu_io_opcode),
    .io_acc_a_data_valid(alu_io_acc_a_data_valid),
    .io_acc_a_data_bits_0_0(alu_io_acc_a_data_bits_0_0),
    .io_acc_a_data_bits_0_1(alu_io_acc_a_data_bits_0_1),
    .io_acc_a_data_bits_0_2(alu_io_acc_a_data_bits_0_2),
    .io_acc_a_data_bits_0_3(alu_io_acc_a_data_bits_0_3),
    .io_acc_a_data_bits_0_4(alu_io_acc_a_data_bits_0_4),
    .io_acc_a_data_bits_0_5(alu_io_acc_a_data_bits_0_5),
    .io_acc_a_data_bits_0_6(alu_io_acc_a_data_bits_0_6),
    .io_acc_a_data_bits_0_7(alu_io_acc_a_data_bits_0_7),
    .io_acc_a_data_bits_0_8(alu_io_acc_a_data_bits_0_8),
    .io_acc_a_data_bits_0_9(alu_io_acc_a_data_bits_0_9),
    .io_acc_a_data_bits_0_10(alu_io_acc_a_data_bits_0_10),
    .io_acc_a_data_bits_0_11(alu_io_acc_a_data_bits_0_11),
    .io_acc_a_data_bits_0_12(alu_io_acc_a_data_bits_0_12),
    .io_acc_a_data_bits_0_13(alu_io_acc_a_data_bits_0_13),
    .io_acc_a_data_bits_0_14(alu_io_acc_a_data_bits_0_14),
    .io_acc_a_data_bits_0_15(alu_io_acc_a_data_bits_0_15),
    .io_acc_b_data_valid(alu_io_acc_b_data_valid),
    .io_acc_b_data_bits_0_0(alu_io_acc_b_data_bits_0_0),
    .io_acc_b_data_bits_0_1(alu_io_acc_b_data_bits_0_1),
    .io_acc_b_data_bits_0_2(alu_io_acc_b_data_bits_0_2),
    .io_acc_b_data_bits_0_3(alu_io_acc_b_data_bits_0_3),
    .io_acc_b_data_bits_0_4(alu_io_acc_b_data_bits_0_4),
    .io_acc_b_data_bits_0_5(alu_io_acc_b_data_bits_0_5),
    .io_acc_b_data_bits_0_6(alu_io_acc_b_data_bits_0_6),
    .io_acc_b_data_bits_0_7(alu_io_acc_b_data_bits_0_7),
    .io_acc_b_data_bits_0_8(alu_io_acc_b_data_bits_0_8),
    .io_acc_b_data_bits_0_9(alu_io_acc_b_data_bits_0_9),
    .io_acc_b_data_bits_0_10(alu_io_acc_b_data_bits_0_10),
    .io_acc_b_data_bits_0_11(alu_io_acc_b_data_bits_0_11),
    .io_acc_b_data_bits_0_12(alu_io_acc_b_data_bits_0_12),
    .io_acc_b_data_bits_0_13(alu_io_acc_b_data_bits_0_13),
    .io_acc_b_data_bits_0_14(alu_io_acc_b_data_bits_0_14),
    .io_acc_b_data_bits_0_15(alu_io_acc_b_data_bits_0_15),
    .io_acc_y_data_valid(alu_io_acc_y_data_valid),
    .io_acc_y_data_bits_0_0(alu_io_acc_y_data_bits_0_0),
    .io_acc_y_data_bits_0_1(alu_io_acc_y_data_bits_0_1),
    .io_acc_y_data_bits_0_2(alu_io_acc_y_data_bits_0_2),
    .io_acc_y_data_bits_0_3(alu_io_acc_y_data_bits_0_3),
    .io_acc_y_data_bits_0_4(alu_io_acc_y_data_bits_0_4),
    .io_acc_y_data_bits_0_5(alu_io_acc_y_data_bits_0_5),
    .io_acc_y_data_bits_0_6(alu_io_acc_y_data_bits_0_6),
    .io_acc_y_data_bits_0_7(alu_io_acc_y_data_bits_0_7),
    .io_acc_y_data_bits_0_8(alu_io_acc_y_data_bits_0_8),
    .io_acc_y_data_bits_0_9(alu_io_acc_y_data_bits_0_9),
    .io_acc_y_data_bits_0_10(alu_io_acc_y_data_bits_0_10),
    .io_acc_y_data_bits_0_11(alu_io_acc_y_data_bits_0_11),
    .io_acc_y_data_bits_0_12(alu_io_acc_y_data_bits_0_12),
    .io_acc_y_data_bits_0_13(alu_io_acc_y_data_bits_0_13),
    .io_acc_y_data_bits_0_14(alu_io_acc_y_data_bits_0_14),
    .io_acc_y_data_bits_0_15(alu_io_acc_y_data_bits_0_15),
    .io_out_data_valid(alu_io_out_data_valid),
    .io_out_data_bits_0_0(alu_io_out_data_bits_0_0),
    .io_out_data_bits_0_1(alu_io_out_data_bits_0_1),
    .io_out_data_bits_0_2(alu_io_out_data_bits_0_2),
    .io_out_data_bits_0_3(alu_io_out_data_bits_0_3),
    .io_out_data_bits_0_4(alu_io_out_data_bits_0_4),
    .io_out_data_bits_0_5(alu_io_out_data_bits_0_5),
    .io_out_data_bits_0_6(alu_io_out_data_bits_0_6),
    .io_out_data_bits_0_7(alu_io_out_data_bits_0_7),
    .io_out_data_bits_0_8(alu_io_out_data_bits_0_8),
    .io_out_data_bits_0_9(alu_io_out_data_bits_0_9),
    .io_out_data_bits_0_10(alu_io_out_data_bits_0_10),
    .io_out_data_bits_0_11(alu_io_out_data_bits_0_11),
    .io_out_data_bits_0_12(alu_io_out_data_bits_0_12),
    .io_out_data_bits_0_13(alu_io_out_data_bits_0_13),
    .io_out_data_bits_0_14(alu_io_out_data_bits_0_14),
    .io_out_data_bits_0_15(alu_io_out_data_bits_0_15)
  );
  assign dec_uop_begin = io_inst[20:8]; // @[TensorAlu.scala 120:29:@22677.4]
  assign dec_uop_end = io_inst[34:21]; // @[TensorAlu.scala 120:29:@22679.4]
  assign dec_lp_0 = io_inst[48:35]; // @[TensorAlu.scala 120:29:@22681.4]
  assign dec_lp_1 = io_inst[62:49]; // @[TensorAlu.scala 120:29:@22683.4]
  assign dec_dst_0 = io_inst[74:64]; // @[TensorAlu.scala 120:29:@22687.4]
  assign dec_dst_1 = io_inst[85:75]; // @[TensorAlu.scala 120:29:@22689.4]
  assign dec_src_0 = io_inst[96:86]; // @[TensorAlu.scala 120:29:@22691.4]
  assign dec_src_1 = io_inst[107:97]; // @[TensorAlu.scala 120:29:@22693.4]
  assign dec_alu_op = io_inst[109:108]; // @[TensorAlu.scala 120:29:@22695.4]
  assign dec_alu_use_imm = io_inst[110]; // @[TensorAlu.scala 120:29:@22697.4]
  assign dec_alu_imm = io_inst[126:111]; // @[TensorAlu.scala 120:29:@22699.4]
  assign _T_1440 = state == 3'h5; // @[TensorAlu.scala 132:11:@22712.4]
  assign _T_1441 = _T_1440 & alu_io_out_data_valid; // @[TensorAlu.scala 132:20:@22713.4]
  assign _T_1443 = dec_lp_0 - 14'h1; // @[TensorAlu.scala 134:27:@22714.4]
  assign _T_1444 = $unsigned(_T_1443); // @[TensorAlu.scala 134:27:@22715.4]
  assign _T_1445 = _T_1444[13:0]; // @[TensorAlu.scala 134:27:@22716.4]
  assign _T_1446 = cnt_o == _T_1445; // @[TensorAlu.scala 134:14:@22717.4]
  assign _T_1447 = _T_1441 & _T_1446; // @[TensorAlu.scala 133:29:@22718.4]
  assign _T_1449 = dec_lp_1 - 14'h1; // @[TensorAlu.scala 135:27:@22719.4]
  assign _T_1450 = $unsigned(_T_1449); // @[TensorAlu.scala 135:27:@22720.4]
  assign _T_1451 = _T_1450[13:0]; // @[TensorAlu.scala 135:27:@22721.4]
  assign _T_1452 = cnt_i == _T_1451; // @[TensorAlu.scala 135:14:@22722.4]
  assign _T_1453 = _T_1447 & _T_1452; // @[TensorAlu.scala 134:34:@22723.4]
  assign _T_1455 = dec_uop_end - 14'h1; // @[TensorAlu.scala 136:28:@22724.4]
  assign _T_1456 = $unsigned(_T_1455); // @[TensorAlu.scala 136:28:@22725.4]
  assign _T_1457 = _T_1456[13:0]; // @[TensorAlu.scala 136:28:@22726.4]
  assign _T_1458 = uop_idx == _T_1457; // @[TensorAlu.scala 136:16:@22727.4]
  assign _T_1459 = 3'h0 == state; // @[Conditional.scala 37:30:@22729.4]
  assign _GEN_0 = io_start ? 3'h1 : state; // @[TensorAlu.scala 140:22:@22731.6]
  assign _T_1460 = 3'h1 == state; // @[Conditional.scala 37:30:@22736.6]
  assign _T_1461 = 3'h2 == state; // @[Conditional.scala 37:30:@22741.8]
  assign _T_1462 = 3'h3 == state; // @[Conditional.scala 37:30:@22746.10]
  assign _T_1463 = 3'h4 == state; // @[Conditional.scala 37:30:@22751.12]
  assign _T_1464 = 3'h5 == state; // @[Conditional.scala 37:30:@22756.14]
  assign _T_1475 = _T_1446 & _T_1452; // @[TensorAlu.scala 159:38:@22767.18]
  assign _T_1481 = _T_1475 & _T_1458; // @[TensorAlu.scala 160:40:@22772.18]
  assign _GEN_1 = _T_1481 ? 3'h0 : 3'h1; // @[TensorAlu.scala 161:42:@22773.18]
  assign _GEN_2 = alu_io_out_data_valid ? _GEN_1 : state; // @[TensorAlu.scala 157:35:@22758.16]
  assign _GEN_3 = _T_1464 ? _GEN_2 : state; // @[Conditional.scala 39:67:@22757.14]
  assign _GEN_4 = _T_1463 ? 3'h5 : _GEN_3; // @[Conditional.scala 39:67:@22752.12]
  assign _GEN_5 = _T_1462 ? 3'h4 : _GEN_4; // @[Conditional.scala 39:67:@22747.10]
  assign _GEN_6 = _T_1461 ? 3'h3 : _GEN_5; // @[Conditional.scala 39:67:@22742.8]
  assign _GEN_7 = _T_1460 ? 3'h2 : _GEN_6; // @[Conditional.scala 39:67:@22737.6]
  assign _GEN_8 = _T_1459 ? _GEN_0 : _GEN_7; // @[Conditional.scala 40:58:@22730.4]
  assign _T_1482 = state == 3'h0; // @[TensorAlu.scala 171:11:@22781.4]
  assign _T_1490 = _T_1441 & _T_1458; // @[TensorAlu.scala 173:31:@22788.4]
  assign _T_1491 = _T_1482 | _T_1490; // @[TensorAlu.scala 171:21:@22789.4]
  assign _T_1495 = uop_idx + 14'h1; // @[TensorAlu.scala 177:24:@22797.8]
  assign _T_1496 = uop_idx + 14'h1; // @[TensorAlu.scala 177:24:@22798.8]
  assign _GEN_9 = _T_1441 ? _T_1496 : uop_idx; // @[TensorAlu.scala 176:55:@22796.6]
  assign _T_1514 = _T_1490 & _T_1452; // @[TensorAlu.scala 187:33:@22819.6]
  assign _T_1516 = cnt_o + 14'h1; // @[TensorAlu.scala 189:20:@22821.8]
  assign _T_1517 = cnt_o + 14'h1; // @[TensorAlu.scala 189:20:@22822.8]
  assign _GEN_28 = {{3'd0}, dec_dst_0}; // @[TensorAlu.scala 190:20:@22824.8]
  assign _T_1518 = dst_o + _GEN_28; // @[TensorAlu.scala 190:20:@22824.8]
  assign _T_1519 = dst_o + _GEN_28; // @[TensorAlu.scala 190:20:@22825.8]
  assign _GEN_29 = {{3'd0}, dec_src_0}; // @[TensorAlu.scala 191:20:@22827.8]
  assign _T_1520 = src_o + _GEN_29; // @[TensorAlu.scala 191:20:@22827.8]
  assign _T_1521 = src_o + _GEN_29; // @[TensorAlu.scala 191:20:@22828.8]
  assign _GEN_11 = _T_1514 ? _T_1517 : cnt_o; // @[TensorAlu.scala 188:33:@22820.6]
  assign _GEN_12 = _T_1514 ? _T_1519 : dst_o; // @[TensorAlu.scala 188:33:@22820.6]
  assign _GEN_13 = _T_1514 ? _T_1521 : src_o; // @[TensorAlu.scala 188:33:@22820.6]
  assign _T_1526 = state == 3'h1; // @[TensorAlu.scala 198:20:@22838.6]
  assign _T_1527 = cnt_i == dec_lp_1; // @[TensorAlu.scala 198:42:@22839.6]
  assign _T_1528 = _T_1526 & _T_1527; // @[TensorAlu.scala 198:33:@22840.6]
  assign _T_1539 = cnt_i + 14'h1; // @[TensorAlu.scala 203:20:@22855.10]
  assign _T_1540 = cnt_i + 14'h1; // @[TensorAlu.scala 203:20:@22856.10]
  assign _GEN_30 = {{3'd0}, dec_dst_1}; // @[TensorAlu.scala 204:20:@22858.10]
  assign _T_1541 = dst_i + _GEN_30; // @[TensorAlu.scala 204:20:@22858.10]
  assign _T_1542 = dst_i + _GEN_30; // @[TensorAlu.scala 204:20:@22859.10]
  assign _GEN_31 = {{3'd0}, dec_src_1}; // @[TensorAlu.scala 205:20:@22861.10]
  assign _T_1543 = src_i + _GEN_31; // @[TensorAlu.scala 205:20:@22861.10]
  assign _T_1544 = src_i + _GEN_31; // @[TensorAlu.scala 205:20:@22862.10]
  assign _GEN_17 = _T_1490 ? _T_1540 : cnt_i; // @[TensorAlu.scala 202:84:@22854.8]
  assign _GEN_18 = _T_1490 ? _T_1542 : dst_i; // @[TensorAlu.scala 202:84:@22854.8]
  assign _GEN_19 = _T_1490 ? _T_1544 : src_i; // @[TensorAlu.scala 202:84:@22854.8]
  assign _GEN_20 = _T_1528 ? 14'h0 : _GEN_17; // @[TensorAlu.scala 198:56:@22841.6]
  assign _GEN_21 = _T_1528 ? dst_o : _GEN_18; // @[TensorAlu.scala 198:56:@22841.6]
  assign _GEN_22 = _T_1528 ? src_o : _GEN_19; // @[TensorAlu.scala 198:56:@22841.6]
  assign _T_1545 = state == 3'h2; // @[TensorAlu.scala 208:14:@22865.4]
  assign _T_1546 = _T_1545 & io_uop_data_valid; // @[TensorAlu.scala 208:30:@22866.4]
  assign _GEN_32 = {{3'd0}, io_uop_data_bits_u0}; // @[TensorAlu.scala 209:36:@22868.6]
  assign _T_1547 = _GEN_32 + dst_i; // @[TensorAlu.scala 209:36:@22868.6]
  assign _T_1548 = _GEN_32 + dst_i; // @[TensorAlu.scala 209:36:@22869.6]
  assign _GEN_33 = {{3'd0}, io_uop_data_bits_u1}; // @[TensorAlu.scala 210:36:@22871.6]
  assign _T_1549 = _GEN_33 + src_i; // @[TensorAlu.scala 210:36:@22871.6]
  assign _T_1550 = _GEN_33 + src_i; // @[TensorAlu.scala 210:36:@22872.6]
  assign _T_1552 = state == 3'h3; // @[TensorAlu.scala 218:32:@22878.4]
  assign _T_1553 = state == 3'h4; // @[TensorAlu.scala 218:58:@22879.4]
  assign _T_1554 = ~ dec_alu_use_imm; // @[TensorAlu.scala 218:77:@22880.4]
  assign _T_1555 = _T_1553 & _T_1554; // @[TensorAlu.scala 218:75:@22881.4]
  assign _T_1558 = _T_1552 ? uop_dst : uop_src; // @[TensorAlu.scala 219:28:@22885.4]
  assign _T_1863 = dec_alu_imm[15]; // @[TensorAlu.scala 226:27:@22890.4]
  assign _T_1866 = {16'hffff,dec_alu_imm}; // @[Cat.scala 30:58:@22892.4]
  assign tensorImm_data_bits_0_0 = _T_1863 ? _T_1866 : {{16'd0}, dec_alu_imm}; // @[TensorAlu.scala 226:15:@22893.4]
  assign _GEN_34 = {{1'd0}, dec_alu_op}; // @[TensorAlu.scala 232:26:@22970.4]
  assign isSHR = _GEN_34 == 3'h3; // @[TensorAlu.scala 232:26:@22970.4]
  assign neg_shift = isSHR & _T_1863; // @[TensorAlu.scala 233:25:@22972.4]
  assign _T_1945 = neg_shift ? 2'h0 : dec_alu_op; // @[TensorAlu.scala 234:40:@22973.4]
  assign _T_1949 = io_acc_rd_data_valid & _T_1440; // @[TensorAlu.scala 240:26:@22996.4]
  assign io_done = _T_1453 & _T_1458; // @[TensorAlu.scala 256:11:@23054.4]
  assign io_uop_idx_valid = state == 3'h1; // @[TensorAlu.scala 214:20:@22876.4]
  assign io_uop_idx_bits = uop_idx[10:0]; // @[TensorAlu.scala 215:19:@22877.4]
  assign io_acc_rd_idx_valid = _T_1552 | _T_1555; // @[TensorAlu.scala 218:23:@22883.4]
  assign io_acc_rd_idx_bits = _T_1558[10:0]; // @[TensorAlu.scala 219:22:@22886.4]
  assign io_acc_wr_valid = alu_io_acc_y_data_valid; // @[TensorAlu.scala 246:19:@23016.4]
  assign io_acc_wr_bits_idx = uop_dst[10:0]; // @[TensorAlu.scala 247:22:@23017.4]
  assign io_acc_wr_bits_data_0_0 = alu_io_acc_y_data_bits_0_0; // @[TensorAlu.scala 248:23:@23018.4]
  assign io_acc_wr_bits_data_0_1 = alu_io_acc_y_data_bits_0_1; // @[TensorAlu.scala 248:23:@23019.4]
  assign io_acc_wr_bits_data_0_2 = alu_io_acc_y_data_bits_0_2; // @[TensorAlu.scala 248:23:@23020.4]
  assign io_acc_wr_bits_data_0_3 = alu_io_acc_y_data_bits_0_3; // @[TensorAlu.scala 248:23:@23021.4]
  assign io_acc_wr_bits_data_0_4 = alu_io_acc_y_data_bits_0_4; // @[TensorAlu.scala 248:23:@23022.4]
  assign io_acc_wr_bits_data_0_5 = alu_io_acc_y_data_bits_0_5; // @[TensorAlu.scala 248:23:@23023.4]
  assign io_acc_wr_bits_data_0_6 = alu_io_acc_y_data_bits_0_6; // @[TensorAlu.scala 248:23:@23024.4]
  assign io_acc_wr_bits_data_0_7 = alu_io_acc_y_data_bits_0_7; // @[TensorAlu.scala 248:23:@23025.4]
  assign io_acc_wr_bits_data_0_8 = alu_io_acc_y_data_bits_0_8; // @[TensorAlu.scala 248:23:@23026.4]
  assign io_acc_wr_bits_data_0_9 = alu_io_acc_y_data_bits_0_9; // @[TensorAlu.scala 248:23:@23027.4]
  assign io_acc_wr_bits_data_0_10 = alu_io_acc_y_data_bits_0_10; // @[TensorAlu.scala 248:23:@23028.4]
  assign io_acc_wr_bits_data_0_11 = alu_io_acc_y_data_bits_0_11; // @[TensorAlu.scala 248:23:@23029.4]
  assign io_acc_wr_bits_data_0_12 = alu_io_acc_y_data_bits_0_12; // @[TensorAlu.scala 248:23:@23030.4]
  assign io_acc_wr_bits_data_0_13 = alu_io_acc_y_data_bits_0_13; // @[TensorAlu.scala 248:23:@23031.4]
  assign io_acc_wr_bits_data_0_14 = alu_io_acc_y_data_bits_0_14; // @[TensorAlu.scala 248:23:@23032.4]
  assign io_acc_wr_bits_data_0_15 = alu_io_acc_y_data_bits_0_15; // @[TensorAlu.scala 248:23:@23033.4]
  assign io_out_wr_valid = alu_io_out_data_valid; // @[TensorAlu.scala 251:19:@23034.4]
  assign io_out_wr_bits_idx = uop_dst[10:0]; // @[TensorAlu.scala 252:22:@23035.4]
  assign io_out_wr_bits_data_0_0 = alu_io_out_data_bits_0_0; // @[TensorAlu.scala 253:23:@23036.4]
  assign io_out_wr_bits_data_0_1 = alu_io_out_data_bits_0_1; // @[TensorAlu.scala 253:23:@23037.4]
  assign io_out_wr_bits_data_0_2 = alu_io_out_data_bits_0_2; // @[TensorAlu.scala 253:23:@23038.4]
  assign io_out_wr_bits_data_0_3 = alu_io_out_data_bits_0_3; // @[TensorAlu.scala 253:23:@23039.4]
  assign io_out_wr_bits_data_0_4 = alu_io_out_data_bits_0_4; // @[TensorAlu.scala 253:23:@23040.4]
  assign io_out_wr_bits_data_0_5 = alu_io_out_data_bits_0_5; // @[TensorAlu.scala 253:23:@23041.4]
  assign io_out_wr_bits_data_0_6 = alu_io_out_data_bits_0_6; // @[TensorAlu.scala 253:23:@23042.4]
  assign io_out_wr_bits_data_0_7 = alu_io_out_data_bits_0_7; // @[TensorAlu.scala 253:23:@23043.4]
  assign io_out_wr_bits_data_0_8 = alu_io_out_data_bits_0_8; // @[TensorAlu.scala 253:23:@23044.4]
  assign io_out_wr_bits_data_0_9 = alu_io_out_data_bits_0_9; // @[TensorAlu.scala 253:23:@23045.4]
  assign io_out_wr_bits_data_0_10 = alu_io_out_data_bits_0_10; // @[TensorAlu.scala 253:23:@23046.4]
  assign io_out_wr_bits_data_0_11 = alu_io_out_data_bits_0_11; // @[TensorAlu.scala 253:23:@23047.4]
  assign io_out_wr_bits_data_0_12 = alu_io_out_data_bits_0_12; // @[TensorAlu.scala 253:23:@23048.4]
  assign io_out_wr_bits_data_0_13 = alu_io_out_data_bits_0_13; // @[TensorAlu.scala 253:23:@23049.4]
  assign io_out_wr_bits_data_0_14 = alu_io_out_data_bits_0_14; // @[TensorAlu.scala 253:23:@23050.4]
  assign io_out_wr_bits_data_0_15 = alu_io_out_data_bits_0_15; // @[TensorAlu.scala 253:23:@23051.4]
  assign alu_clock = clock; // @[:@22660.4]
  assign alu_io_opcode = {neg_shift,_T_1945}; // @[TensorAlu.scala 235:17:@22975.4]
  assign alu_io_acc_a_data_valid = io_acc_rd_data_valid & _T_1553; // @[TensorAlu.scala 236:27:@22978.4]
  assign alu_io_acc_a_data_bits_0_0 = io_acc_rd_data_bits_0_0; // @[TensorAlu.scala 237:26:@22979.4]
  assign alu_io_acc_a_data_bits_0_1 = io_acc_rd_data_bits_0_1; // @[TensorAlu.scala 237:26:@22980.4]
  assign alu_io_acc_a_data_bits_0_2 = io_acc_rd_data_bits_0_2; // @[TensorAlu.scala 237:26:@22981.4]
  assign alu_io_acc_a_data_bits_0_3 = io_acc_rd_data_bits_0_3; // @[TensorAlu.scala 237:26:@22982.4]
  assign alu_io_acc_a_data_bits_0_4 = io_acc_rd_data_bits_0_4; // @[TensorAlu.scala 237:26:@22983.4]
  assign alu_io_acc_a_data_bits_0_5 = io_acc_rd_data_bits_0_5; // @[TensorAlu.scala 237:26:@22984.4]
  assign alu_io_acc_a_data_bits_0_6 = io_acc_rd_data_bits_0_6; // @[TensorAlu.scala 237:26:@22985.4]
  assign alu_io_acc_a_data_bits_0_7 = io_acc_rd_data_bits_0_7; // @[TensorAlu.scala 237:26:@22986.4]
  assign alu_io_acc_a_data_bits_0_8 = io_acc_rd_data_bits_0_8; // @[TensorAlu.scala 237:26:@22987.4]
  assign alu_io_acc_a_data_bits_0_9 = io_acc_rd_data_bits_0_9; // @[TensorAlu.scala 237:26:@22988.4]
  assign alu_io_acc_a_data_bits_0_10 = io_acc_rd_data_bits_0_10; // @[TensorAlu.scala 237:26:@22989.4]
  assign alu_io_acc_a_data_bits_0_11 = io_acc_rd_data_bits_0_11; // @[TensorAlu.scala 237:26:@22990.4]
  assign alu_io_acc_a_data_bits_0_12 = io_acc_rd_data_bits_0_12; // @[TensorAlu.scala 237:26:@22991.4]
  assign alu_io_acc_a_data_bits_0_13 = io_acc_rd_data_bits_0_13; // @[TensorAlu.scala 237:26:@22992.4]
  assign alu_io_acc_a_data_bits_0_14 = io_acc_rd_data_bits_0_14; // @[TensorAlu.scala 237:26:@22993.4]
  assign alu_io_acc_a_data_bits_0_15 = io_acc_rd_data_bits_0_15; // @[TensorAlu.scala 237:26:@22994.4]
  assign alu_io_acc_b_data_valid = dec_alu_use_imm ? _T_1553 : _T_1949; // @[TensorAlu.scala 238:27:@22998.4]
  assign alu_io_acc_b_data_bits_0_0 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_0; // @[TensorAlu.scala 241:26:@23000.4]
  assign alu_io_acc_b_data_bits_0_1 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_1; // @[TensorAlu.scala 241:26:@23001.4]
  assign alu_io_acc_b_data_bits_0_2 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_2; // @[TensorAlu.scala 241:26:@23002.4]
  assign alu_io_acc_b_data_bits_0_3 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_3; // @[TensorAlu.scala 241:26:@23003.4]
  assign alu_io_acc_b_data_bits_0_4 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_4; // @[TensorAlu.scala 241:26:@23004.4]
  assign alu_io_acc_b_data_bits_0_5 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_5; // @[TensorAlu.scala 241:26:@23005.4]
  assign alu_io_acc_b_data_bits_0_6 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_6; // @[TensorAlu.scala 241:26:@23006.4]
  assign alu_io_acc_b_data_bits_0_7 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_7; // @[TensorAlu.scala 241:26:@23007.4]
  assign alu_io_acc_b_data_bits_0_8 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_8; // @[TensorAlu.scala 241:26:@23008.4]
  assign alu_io_acc_b_data_bits_0_9 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_9; // @[TensorAlu.scala 241:26:@23009.4]
  assign alu_io_acc_b_data_bits_0_10 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_10; // @[TensorAlu.scala 241:26:@23010.4]
  assign alu_io_acc_b_data_bits_0_11 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_11; // @[TensorAlu.scala 241:26:@23011.4]
  assign alu_io_acc_b_data_bits_0_12 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_12; // @[TensorAlu.scala 241:26:@23012.4]
  assign alu_io_acc_b_data_bits_0_13 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_13; // @[TensorAlu.scala 241:26:@23013.4]
  assign alu_io_acc_b_data_bits_0_14 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_14; // @[TensorAlu.scala 241:26:@23014.4]
  assign alu_io_acc_b_data_bits_0_15 = dec_alu_use_imm ? tensorImm_data_bits_0_0 : io_acc_rd_data_bits_0_15; // @[TensorAlu.scala 241:26:@23015.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  uop_idx = _RAND_1[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  uop_dst = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  uop_src = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cnt_o = _RAND_4[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  dst_o = _RAND_5[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  src_o = _RAND_6[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  cnt_i = _RAND_7[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  dst_i = _RAND_8[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  src_i = _RAND_9[13:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_1459) begin
        if (io_start) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_1460) begin
          state <= 3'h2;
        end else begin
          if (_T_1461) begin
            state <= 3'h3;
          end else begin
            if (_T_1462) begin
              state <= 3'h4;
            end else begin
              if (_T_1463) begin
                state <= 3'h5;
              end else begin
                if (_T_1464) begin
                  if (alu_io_out_data_valid) begin
                    if (_T_1481) begin
                      state <= 3'h0;
                    end else begin
                      state <= 3'h1;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_1491) begin
      uop_idx <= {{1'd0}, dec_uop_begin};
    end else begin
      if (_T_1441) begin
        uop_idx <= _T_1496;
      end
    end
    if (_T_1546) begin
      uop_dst <= _T_1548;
    end
    if (_T_1546) begin
      uop_src <= _T_1550;
    end
    if (_T_1482) begin
      cnt_o <= 14'h0;
    end else begin
      if (_T_1514) begin
        cnt_o <= _T_1517;
      end
    end
    if (_T_1482) begin
      dst_o <= 14'h0;
    end else begin
      if (_T_1514) begin
        dst_o <= _T_1519;
      end
    end
    if (_T_1482) begin
      src_o <= 14'h0;
    end else begin
      if (_T_1514) begin
        src_o <= _T_1521;
      end
    end
    if (_T_1482) begin
      cnt_i <= 14'h0;
    end else begin
      if (_T_1528) begin
        cnt_i <= 14'h0;
      end else begin
        if (_T_1490) begin
          cnt_i <= _T_1540;
        end
      end
    end
    if (_T_1482) begin
      dst_i <= 14'h0;
    end else begin
      if (_T_1528) begin
        dst_i <= dst_o;
      end else begin
        if (_T_1490) begin
          dst_i <= _T_1542;
        end
      end
    end
    if (_T_1482) begin
      src_i <= 14'h0;
    end else begin
      if (_T_1528) begin
        src_i <= src_o;
      end else begin
        if (_T_1490) begin
          src_i <= _T_1544;
        end
      end
    end
  end
endmodule
module ComputeDecode( // @[:@23107.2]
  input  [127:0] io_inst, // @[:@23110.4]
  output         io_push_next, // @[:@23110.4]
  output         io_push_prev, // @[:@23110.4]
  output         io_pop_next, // @[:@23110.4]
  output         io_pop_prev, // @[:@23110.4]
  output         io_isLoadAcc, // @[:@23110.4]
  output         io_isLoadUop, // @[:@23110.4]
  output         io_isSync, // @[:@23110.4]
  output         io_isAlu, // @[:@23110.4]
  output         io_isGemm, // @[:@23110.4]
  output         io_isFinish // @[:@23110.4]
);
  wire [15:0] dec_xsize; // @[Decode.scala 200:29:@23135.4]
  wire [127:0] _T_49; // @[Decode.scala 205:27:@23151.4]
  wire  _T_50; // @[Decode.scala 205:27:@23152.4]
  wire  _T_52; // @[Decode.scala 205:48:@23153.4]
  wire  _T_57; // @[Decode.scala 206:27:@23157.4]
  wire  _T_69; // @[Decode.scala 207:34:@23165.4]
  wire  _T_71; // @[Decode.scala 207:66:@23166.4]
  wire [127:0] _T_75; // @[Decode.scala 208:23:@23169.4]
  wire  _T_76; // @[Decode.scala 208:23:@23170.4]
  wire  _T_80; // @[Decode.scala 208:42:@23172.4]
  wire  _T_81; // @[Decode.scala 208:32:@23173.4]
  wire  _T_85; // @[Decode.scala 208:61:@23175.4]
  wire  _T_86; // @[Decode.scala 208:51:@23176.4]
  wire  _T_90; // @[Decode.scala 208:80:@23178.4]
  wire [127:0] _T_94; // @[Decode.scala 209:24:@23181.4]
  assign dec_xsize = io_inst[95:80]; // @[Decode.scala 200:29:@23135.4]
  assign _T_49 = io_inst & 128'h187; // @[Decode.scala 205:27:@23151.4]
  assign _T_50 = 128'h180 == _T_49; // @[Decode.scala 205:27:@23152.4]
  assign _T_52 = dec_xsize != 16'h0; // @[Decode.scala 205:48:@23153.4]
  assign _T_57 = 128'h0 == _T_49; // @[Decode.scala 206:27:@23157.4]
  assign _T_69 = _T_50 | _T_57; // @[Decode.scala 207:34:@23165.4]
  assign _T_71 = dec_xsize == 16'h0; // @[Decode.scala 207:66:@23166.4]
  assign _T_75 = io_inst & 128'h3000000000000000000000000007; // @[Decode.scala 208:23:@23169.4]
  assign _T_76 = 128'h4 == _T_75; // @[Decode.scala 208:23:@23170.4]
  assign _T_80 = 128'h1000000000000000000000000004 == _T_75; // @[Decode.scala 208:42:@23172.4]
  assign _T_81 = _T_76 | _T_80; // @[Decode.scala 208:32:@23173.4]
  assign _T_85 = 128'h2000000000000000000000000004 == _T_75; // @[Decode.scala 208:61:@23175.4]
  assign _T_86 = _T_81 | _T_85; // @[Decode.scala 208:51:@23176.4]
  assign _T_90 = 128'h3000000000000000000000000004 == _T_75; // @[Decode.scala 208:80:@23178.4]
  assign _T_94 = io_inst & 128'h7; // @[Decode.scala 209:24:@23181.4]
  assign io_push_next = io_inst[6]; // @[Decode.scala 201:16:@23147.4]
  assign io_push_prev = io_inst[5]; // @[Decode.scala 202:16:@23148.4]
  assign io_pop_next = io_inst[4]; // @[Decode.scala 203:15:@23149.4]
  assign io_pop_prev = io_inst[3]; // @[Decode.scala 204:15:@23150.4]
  assign io_isLoadAcc = _T_50 & _T_52; // @[Decode.scala 205:16:@23155.4]
  assign io_isLoadUop = _T_57 & _T_52; // @[Decode.scala 206:16:@23160.4]
  assign io_isSync = _T_69 & _T_71; // @[Decode.scala 207:13:@23168.4]
  assign io_isAlu = _T_86 | _T_90; // @[Decode.scala 208:12:@23180.4]
  assign io_isGemm = 128'h2 == _T_94; // @[Decode.scala 209:13:@23183.4]
  assign io_isFinish = 128'h3 == _T_94; // @[Decode.scala 210:15:@23186.4]
endmodule
module Compute( // @[:@23188.2]
  input          clock, // @[:@23189.4]
  input          reset, // @[:@23190.4]
  input          io_i_post_0, // @[:@23191.4]
  input          io_i_post_1, // @[:@23191.4]
  output         io_o_post_0, // @[:@23191.4]
  output         io_o_post_1, // @[:@23191.4]
  output         io_inst_ready, // @[:@23191.4]
  input          io_inst_valid, // @[:@23191.4]
  input  [127:0] io_inst_bits, // @[:@23191.4]
  input  [31:0]  io_uop_baddr, // @[:@23191.4]
  input  [31:0]  io_acc_baddr, // @[:@23191.4]
  input          io_vme_rd_0_cmd_ready, // @[:@23191.4]
  output         io_vme_rd_0_cmd_valid, // @[:@23191.4]
  output [31:0]  io_vme_rd_0_cmd_bits_addr, // @[:@23191.4]
  output [7:0]   io_vme_rd_0_cmd_bits_len, // @[:@23191.4]
  output         io_vme_rd_0_data_ready, // @[:@23191.4]
  input          io_vme_rd_0_data_valid, // @[:@23191.4]
  input  [63:0]  io_vme_rd_0_data_bits, // @[:@23191.4]
  input          io_vme_rd_1_cmd_ready, // @[:@23191.4]
  output         io_vme_rd_1_cmd_valid, // @[:@23191.4]
  output [31:0]  io_vme_rd_1_cmd_bits_addr, // @[:@23191.4]
  output [7:0]   io_vme_rd_1_cmd_bits_len, // @[:@23191.4]
  output         io_vme_rd_1_data_ready, // @[:@23191.4]
  input          io_vme_rd_1_data_valid, // @[:@23191.4]
  input  [63:0]  io_vme_rd_1_data_bits, // @[:@23191.4]
  output         io_inp_rd_idx_valid, // @[:@23191.4]
  output [10:0]  io_inp_rd_idx_bits, // @[:@23191.4]
  input          io_inp_rd_data_valid, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_0, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_1, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_2, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_3, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_4, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_5, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_6, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_7, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_8, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_9, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_10, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_11, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_12, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_13, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_14, // @[:@23191.4]
  input  [7:0]   io_inp_rd_data_bits_0_15, // @[:@23191.4]
  output         io_wgt_rd_idx_valid, // @[:@23191.4]
  output [9:0]   io_wgt_rd_idx_bits, // @[:@23191.4]
  input          io_wgt_rd_data_valid, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_0_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_1_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_2_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_3_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_4_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_5_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_6_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_7_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_8_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_9_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_10_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_11_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_12_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_13_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_14_15, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_0, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_1, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_2, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_3, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_4, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_5, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_6, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_7, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_8, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_9, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_10, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_11, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_12, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_13, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_14, // @[:@23191.4]
  input  [7:0]   io_wgt_rd_data_bits_15_15, // @[:@23191.4]
  output         io_out_wr_valid, // @[:@23191.4]
  output [10:0]  io_out_wr_bits_idx, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_0, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_1, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_2, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_3, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_4, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_5, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_6, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_7, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_8, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_9, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_10, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_11, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_12, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_13, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_14, // @[:@23191.4]
  output [7:0]   io_out_wr_bits_data_0_15, // @[:@23191.4]
  output         io_finish, // @[:@23191.4]
  output         io_acc_wr_event // @[:@23191.4]
);
  wire  s_0_clock; // @[Compute.scala 54:11:@23194.4]
  wire  s_0_reset; // @[Compute.scala 54:11:@23194.4]
  wire  s_0_io_spost; // @[Compute.scala 54:11:@23194.4]
  wire  s_0_io_swait; // @[Compute.scala 54:11:@23194.4]
  wire  s_0_io_sready; // @[Compute.scala 54:11:@23194.4]
  wire  s_1_clock; // @[Compute.scala 54:11:@23197.4]
  wire  s_1_reset; // @[Compute.scala 54:11:@23197.4]
  wire  s_1_io_spost; // @[Compute.scala 54:11:@23197.4]
  wire  s_1_io_swait; // @[Compute.scala 54:11:@23197.4]
  wire  s_1_io_sready; // @[Compute.scala 54:11:@23197.4]
  wire  loadUop_clock; // @[Compute.scala 56:23:@23200.4]
  wire  loadUop_reset; // @[Compute.scala 56:23:@23200.4]
  wire  loadUop_io_start; // @[Compute.scala 56:23:@23200.4]
  wire  loadUop_io_done; // @[Compute.scala 56:23:@23200.4]
  wire [127:0] loadUop_io_inst; // @[Compute.scala 56:23:@23200.4]
  wire [31:0] loadUop_io_baddr; // @[Compute.scala 56:23:@23200.4]
  wire  loadUop_io_vme_rd_cmd_ready; // @[Compute.scala 56:23:@23200.4]
  wire  loadUop_io_vme_rd_cmd_valid; // @[Compute.scala 56:23:@23200.4]
  wire [31:0] loadUop_io_vme_rd_cmd_bits_addr; // @[Compute.scala 56:23:@23200.4]
  wire [7:0] loadUop_io_vme_rd_cmd_bits_len; // @[Compute.scala 56:23:@23200.4]
  wire  loadUop_io_vme_rd_data_ready; // @[Compute.scala 56:23:@23200.4]
  wire  loadUop_io_vme_rd_data_valid; // @[Compute.scala 56:23:@23200.4]
  wire [63:0] loadUop_io_vme_rd_data_bits; // @[Compute.scala 56:23:@23200.4]
  wire  loadUop_io_uop_idx_valid; // @[Compute.scala 56:23:@23200.4]
  wire [10:0] loadUop_io_uop_idx_bits; // @[Compute.scala 56:23:@23200.4]
  wire  loadUop_io_uop_data_valid; // @[Compute.scala 56:23:@23200.4]
  wire [9:0] loadUop_io_uop_data_bits_u2; // @[Compute.scala 56:23:@23200.4]
  wire [10:0] loadUop_io_uop_data_bits_u1; // @[Compute.scala 56:23:@23200.4]
  wire [10:0] loadUop_io_uop_data_bits_u0; // @[Compute.scala 56:23:@23200.4]
  wire  tensorAcc_clock; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_reset; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_io_start; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_io_done; // @[Compute.scala 57:25:@23203.4]
  wire [127:0] tensorAcc_io_inst; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_baddr; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_io_vme_rd_cmd_ready; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_io_vme_rd_cmd_valid; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_vme_rd_cmd_bits_addr; // @[Compute.scala 57:25:@23203.4]
  wire [7:0] tensorAcc_io_vme_rd_cmd_bits_len; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_io_vme_rd_data_ready; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_io_vme_rd_data_valid; // @[Compute.scala 57:25:@23203.4]
  wire [63:0] tensorAcc_io_vme_rd_data_bits; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_io_tensor_rd_idx_valid; // @[Compute.scala 57:25:@23203.4]
  wire [10:0] tensorAcc_io_tensor_rd_idx_bits; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_io_tensor_rd_data_valid; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_0; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_1; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_2; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_3; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_4; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_5; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_6; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_7; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_8; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_9; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_10; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_11; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_12; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_13; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_14; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_rd_data_bits_0_15; // @[Compute.scala 57:25:@23203.4]
  wire  tensorAcc_io_tensor_wr_valid; // @[Compute.scala 57:25:@23203.4]
  wire [10:0] tensorAcc_io_tensor_wr_bits_idx; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_0; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_1; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_2; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_3; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_4; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_5; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_6; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_7; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_8; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_9; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_10; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_11; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_12; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_13; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_14; // @[Compute.scala 57:25:@23203.4]
  wire [31:0] tensorAcc_io_tensor_wr_bits_data_0_15; // @[Compute.scala 57:25:@23203.4]
  wire  tensorGemm_clock; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_reset; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_start; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_done; // @[Compute.scala 58:26:@23206.4]
  wire [127:0] tensorGemm_io_inst; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_uop_idx_valid; // @[Compute.scala 58:26:@23206.4]
  wire [10:0] tensorGemm_io_uop_idx_bits; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_uop_data_valid; // @[Compute.scala 58:26:@23206.4]
  wire [9:0] tensorGemm_io_uop_data_bits_u2; // @[Compute.scala 58:26:@23206.4]
  wire [10:0] tensorGemm_io_uop_data_bits_u1; // @[Compute.scala 58:26:@23206.4]
  wire [10:0] tensorGemm_io_uop_data_bits_u0; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_inp_rd_idx_valid; // @[Compute.scala 58:26:@23206.4]
  wire [10:0] tensorGemm_io_inp_rd_idx_bits; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_inp_rd_data_valid; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_inp_rd_data_bits_0_15; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_wgt_rd_idx_valid; // @[Compute.scala 58:26:@23206.4]
  wire [9:0] tensorGemm_io_wgt_rd_idx_bits; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_wgt_rd_data_valid; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_0_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_1_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_2_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_3_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_4_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_5_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_6_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_7_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_8_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_9_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_10_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_11_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_12_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_13_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_14_15; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_wgt_rd_data_bits_15_15; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_acc_rd_idx_valid; // @[Compute.scala 58:26:@23206.4]
  wire [10:0] tensorGemm_io_acc_rd_idx_bits; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_acc_rd_data_valid; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_0; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_1; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_2; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_3; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_4; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_5; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_6; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_7; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_8; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_9; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_10; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_11; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_12; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_13; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_14; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_rd_data_bits_0_15; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_acc_wr_valid; // @[Compute.scala 58:26:@23206.4]
  wire [10:0] tensorGemm_io_acc_wr_bits_idx; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_0; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_1; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_2; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_3; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_4; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_5; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_6; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_7; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_8; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_9; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_10; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_11; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_12; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_13; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_14; // @[Compute.scala 58:26:@23206.4]
  wire [31:0] tensorGemm_io_acc_wr_bits_data_0_15; // @[Compute.scala 58:26:@23206.4]
  wire  tensorGemm_io_out_wr_valid; // @[Compute.scala 58:26:@23206.4]
  wire [10:0] tensorGemm_io_out_wr_bits_idx; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_0; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_1; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_2; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_3; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_4; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_5; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_6; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_7; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_8; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_9; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_10; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_11; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_12; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_13; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_14; // @[Compute.scala 58:26:@23206.4]
  wire [7:0] tensorGemm_io_out_wr_bits_data_0_15; // @[Compute.scala 58:26:@23206.4]
  wire  tensorAlu_clock; // @[Compute.scala 59:25:@23209.4]
  wire  tensorAlu_reset; // @[Compute.scala 59:25:@23209.4]
  wire  tensorAlu_io_start; // @[Compute.scala 59:25:@23209.4]
  wire  tensorAlu_io_done; // @[Compute.scala 59:25:@23209.4]
  wire [127:0] tensorAlu_io_inst; // @[Compute.scala 59:25:@23209.4]
  wire  tensorAlu_io_uop_idx_valid; // @[Compute.scala 59:25:@23209.4]
  wire [10:0] tensorAlu_io_uop_idx_bits; // @[Compute.scala 59:25:@23209.4]
  wire  tensorAlu_io_uop_data_valid; // @[Compute.scala 59:25:@23209.4]
  wire [10:0] tensorAlu_io_uop_data_bits_u1; // @[Compute.scala 59:25:@23209.4]
  wire [10:0] tensorAlu_io_uop_data_bits_u0; // @[Compute.scala 59:25:@23209.4]
  wire  tensorAlu_io_acc_rd_idx_valid; // @[Compute.scala 59:25:@23209.4]
  wire [10:0] tensorAlu_io_acc_rd_idx_bits; // @[Compute.scala 59:25:@23209.4]
  wire  tensorAlu_io_acc_rd_data_valid; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_0; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_1; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_2; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_3; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_4; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_5; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_6; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_7; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_8; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_9; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_10; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_11; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_12; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_13; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_14; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_rd_data_bits_0_15; // @[Compute.scala 59:25:@23209.4]
  wire  tensorAlu_io_acc_wr_valid; // @[Compute.scala 59:25:@23209.4]
  wire [10:0] tensorAlu_io_acc_wr_bits_idx; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_0; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_1; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_2; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_3; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_4; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_5; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_6; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_7; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_8; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_9; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_10; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_11; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_12; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_13; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_14; // @[Compute.scala 59:25:@23209.4]
  wire [31:0] tensorAlu_io_acc_wr_bits_data_0_15; // @[Compute.scala 59:25:@23209.4]
  wire  tensorAlu_io_out_wr_valid; // @[Compute.scala 59:25:@23209.4]
  wire [10:0] tensorAlu_io_out_wr_bits_idx; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_0; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_1; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_2; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_3; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_4; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_5; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_6; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_7; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_8; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_9; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_10; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_11; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_12; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_13; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_14; // @[Compute.scala 59:25:@23209.4]
  wire [7:0] tensorAlu_io_out_wr_bits_data_0_15; // @[Compute.scala 59:25:@23209.4]
  wire  inst_q_clock; // @[Compute.scala 61:22:@23212.4]
  wire  inst_q_reset; // @[Compute.scala 61:22:@23212.4]
  wire  inst_q_io_enq_ready; // @[Compute.scala 61:22:@23212.4]
  wire  inst_q_io_enq_valid; // @[Compute.scala 61:22:@23212.4]
  wire [127:0] inst_q_io_enq_bits; // @[Compute.scala 61:22:@23212.4]
  wire  inst_q_io_deq_ready; // @[Compute.scala 61:22:@23212.4]
  wire  inst_q_io_deq_valid; // @[Compute.scala 61:22:@23212.4]
  wire [127:0] inst_q_io_deq_bits; // @[Compute.scala 61:22:@23212.4]
  wire [127:0] dec_io_inst; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_push_next; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_push_prev; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_pop_next; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_pop_prev; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_isLoadAcc; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_isLoadUop; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_isSync; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_isAlu; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_isGemm; // @[Compute.scala 64:19:@23215.4]
  wire  dec_io_isFinish; // @[Compute.scala 64:19:@23215.4]
  reg [1:0] state; // @[Compute.scala 51:22:@23193.4]
  reg [31:0] _RAND_0;
  wire [4:0] inst_type; // @[Cat.scala 30:58:@23222.4]
  wire  _T_7054; // @[Compute.scala 74:40:@23223.4]
  wire  sprev; // @[Compute.scala 74:35:@23224.4]
  wire  _T_7056; // @[Compute.scala 75:40:@23225.4]
  wire  snext; // @[Compute.scala 75:35:@23226.4]
  wire  start; // @[Compute.scala 76:21:@23227.4]
  wire  _T_7064; // @[Mux.scala 46:19:@23228.4]
  wire  _T_7066; // @[Mux.scala 46:19:@23230.4]
  wire  _T_7067; // @[Mux.scala 46:16:@23231.4]
  wire  _T_7068; // @[Mux.scala 46:19:@23232.4]
  wire  _T_7069; // @[Mux.scala 46:16:@23233.4]
  wire  _T_7070; // @[Mux.scala 46:19:@23234.4]
  wire  _T_7071; // @[Mux.scala 46:16:@23235.4]
  wire  _T_7072; // @[Mux.scala 46:19:@23236.4]
  wire  done; // @[Mux.scala 46:16:@23237.4]
  wire  _T_7073; // @[Conditional.scala 37:30:@23238.4]
  wire  _T_7075; // @[Compute.scala 96:30:@23245.10]
  wire [1:0] _GEN_0; // @[Compute.scala 96:35:@23246.10]
  wire [1:0] _GEN_1; // @[Compute.scala 94:29:@23241.8]
  wire [1:0] _GEN_2; // @[Compute.scala 93:19:@23240.6]
  wire  _T_7076; // @[Conditional.scala 37:30:@23252.6]
  wire  _T_7077; // @[Conditional.scala 37:30:@23257.8]
  wire [1:0] _GEN_3; // @[Compute.scala 105:18:@23259.10]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@23258.8]
  wire [1:0] _GEN_5; // @[Conditional.scala 39:67:@23253.6]
  wire [1:0] _GEN_6; // @[Conditional.scala 40:58:@23239.4]
  wire  _T_7078; // @[Compute.scala 113:33:@23266.4]
  wire  _T_7079; // @[Compute.scala 113:42:@23267.4]
  wire  _T_7080; // @[Compute.scala 113:59:@23268.4]
  wire  _T_7081; // @[Compute.scala 113:50:@23269.4]
  wire  _T_7082; // @[Compute.scala 116:29:@23271.4]
  wire  _T_7083; // @[Compute.scala 116:39:@23272.4]
  Semaphore s_0 ( // @[Compute.scala 54:11:@23194.4]
    .clock(s_0_clock),
    .reset(s_0_reset),
    .io_spost(s_0_io_spost),
    .io_swait(s_0_io_swait),
    .io_sready(s_0_io_sready)
  );
  Semaphore s_1 ( // @[Compute.scala 54:11:@23197.4]
    .clock(s_1_clock),
    .reset(s_1_reset),
    .io_spost(s_1_io_spost),
    .io_swait(s_1_io_swait),
    .io_sready(s_1_io_sready)
  );
  LoadUop loadUop ( // @[Compute.scala 56:23:@23200.4]
    .clock(loadUop_clock),
    .reset(loadUop_reset),
    .io_start(loadUop_io_start),
    .io_done(loadUop_io_done),
    .io_inst(loadUop_io_inst),
    .io_baddr(loadUop_io_baddr),
    .io_vme_rd_cmd_ready(loadUop_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(loadUop_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(loadUop_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(loadUop_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(loadUop_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(loadUop_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(loadUop_io_vme_rd_data_bits),
    .io_uop_idx_valid(loadUop_io_uop_idx_valid),
    .io_uop_idx_bits(loadUop_io_uop_idx_bits),
    .io_uop_data_valid(loadUop_io_uop_data_valid),
    .io_uop_data_bits_u2(loadUop_io_uop_data_bits_u2),
    .io_uop_data_bits_u1(loadUop_io_uop_data_bits_u1),
    .io_uop_data_bits_u0(loadUop_io_uop_data_bits_u0)
  );
  TensorLoad_2 tensorAcc ( // @[Compute.scala 57:25:@23203.4]
    .clock(tensorAcc_clock),
    .reset(tensorAcc_reset),
    .io_start(tensorAcc_io_start),
    .io_done(tensorAcc_io_done),
    .io_inst(tensorAcc_io_inst),
    .io_baddr(tensorAcc_io_baddr),
    .io_vme_rd_cmd_ready(tensorAcc_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorAcc_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorAcc_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorAcc_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(tensorAcc_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorAcc_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(tensorAcc_io_vme_rd_data_bits),
    .io_tensor_rd_idx_valid(tensorAcc_io_tensor_rd_idx_valid),
    .io_tensor_rd_idx_bits(tensorAcc_io_tensor_rd_idx_bits),
    .io_tensor_rd_data_valid(tensorAcc_io_tensor_rd_data_valid),
    .io_tensor_rd_data_bits_0_0(tensorAcc_io_tensor_rd_data_bits_0_0),
    .io_tensor_rd_data_bits_0_1(tensorAcc_io_tensor_rd_data_bits_0_1),
    .io_tensor_rd_data_bits_0_2(tensorAcc_io_tensor_rd_data_bits_0_2),
    .io_tensor_rd_data_bits_0_3(tensorAcc_io_tensor_rd_data_bits_0_3),
    .io_tensor_rd_data_bits_0_4(tensorAcc_io_tensor_rd_data_bits_0_4),
    .io_tensor_rd_data_bits_0_5(tensorAcc_io_tensor_rd_data_bits_0_5),
    .io_tensor_rd_data_bits_0_6(tensorAcc_io_tensor_rd_data_bits_0_6),
    .io_tensor_rd_data_bits_0_7(tensorAcc_io_tensor_rd_data_bits_0_7),
    .io_tensor_rd_data_bits_0_8(tensorAcc_io_tensor_rd_data_bits_0_8),
    .io_tensor_rd_data_bits_0_9(tensorAcc_io_tensor_rd_data_bits_0_9),
    .io_tensor_rd_data_bits_0_10(tensorAcc_io_tensor_rd_data_bits_0_10),
    .io_tensor_rd_data_bits_0_11(tensorAcc_io_tensor_rd_data_bits_0_11),
    .io_tensor_rd_data_bits_0_12(tensorAcc_io_tensor_rd_data_bits_0_12),
    .io_tensor_rd_data_bits_0_13(tensorAcc_io_tensor_rd_data_bits_0_13),
    .io_tensor_rd_data_bits_0_14(tensorAcc_io_tensor_rd_data_bits_0_14),
    .io_tensor_rd_data_bits_0_15(tensorAcc_io_tensor_rd_data_bits_0_15),
    .io_tensor_wr_valid(tensorAcc_io_tensor_wr_valid),
    .io_tensor_wr_bits_idx(tensorAcc_io_tensor_wr_bits_idx),
    .io_tensor_wr_bits_data_0_0(tensorAcc_io_tensor_wr_bits_data_0_0),
    .io_tensor_wr_bits_data_0_1(tensorAcc_io_tensor_wr_bits_data_0_1),
    .io_tensor_wr_bits_data_0_2(tensorAcc_io_tensor_wr_bits_data_0_2),
    .io_tensor_wr_bits_data_0_3(tensorAcc_io_tensor_wr_bits_data_0_3),
    .io_tensor_wr_bits_data_0_4(tensorAcc_io_tensor_wr_bits_data_0_4),
    .io_tensor_wr_bits_data_0_5(tensorAcc_io_tensor_wr_bits_data_0_5),
    .io_tensor_wr_bits_data_0_6(tensorAcc_io_tensor_wr_bits_data_0_6),
    .io_tensor_wr_bits_data_0_7(tensorAcc_io_tensor_wr_bits_data_0_7),
    .io_tensor_wr_bits_data_0_8(tensorAcc_io_tensor_wr_bits_data_0_8),
    .io_tensor_wr_bits_data_0_9(tensorAcc_io_tensor_wr_bits_data_0_9),
    .io_tensor_wr_bits_data_0_10(tensorAcc_io_tensor_wr_bits_data_0_10),
    .io_tensor_wr_bits_data_0_11(tensorAcc_io_tensor_wr_bits_data_0_11),
    .io_tensor_wr_bits_data_0_12(tensorAcc_io_tensor_wr_bits_data_0_12),
    .io_tensor_wr_bits_data_0_13(tensorAcc_io_tensor_wr_bits_data_0_13),
    .io_tensor_wr_bits_data_0_14(tensorAcc_io_tensor_wr_bits_data_0_14),
    .io_tensor_wr_bits_data_0_15(tensorAcc_io_tensor_wr_bits_data_0_15)
  );
  TensorGemm tensorGemm ( // @[Compute.scala 58:26:@23206.4]
    .clock(tensorGemm_clock),
    .reset(tensorGemm_reset),
    .io_start(tensorGemm_io_start),
    .io_done(tensorGemm_io_done),
    .io_inst(tensorGemm_io_inst),
    .io_uop_idx_valid(tensorGemm_io_uop_idx_valid),
    .io_uop_idx_bits(tensorGemm_io_uop_idx_bits),
    .io_uop_data_valid(tensorGemm_io_uop_data_valid),
    .io_uop_data_bits_u2(tensorGemm_io_uop_data_bits_u2),
    .io_uop_data_bits_u1(tensorGemm_io_uop_data_bits_u1),
    .io_uop_data_bits_u0(tensorGemm_io_uop_data_bits_u0),
    .io_inp_rd_idx_valid(tensorGemm_io_inp_rd_idx_valid),
    .io_inp_rd_idx_bits(tensorGemm_io_inp_rd_idx_bits),
    .io_inp_rd_data_valid(tensorGemm_io_inp_rd_data_valid),
    .io_inp_rd_data_bits_0_0(tensorGemm_io_inp_rd_data_bits_0_0),
    .io_inp_rd_data_bits_0_1(tensorGemm_io_inp_rd_data_bits_0_1),
    .io_inp_rd_data_bits_0_2(tensorGemm_io_inp_rd_data_bits_0_2),
    .io_inp_rd_data_bits_0_3(tensorGemm_io_inp_rd_data_bits_0_3),
    .io_inp_rd_data_bits_0_4(tensorGemm_io_inp_rd_data_bits_0_4),
    .io_inp_rd_data_bits_0_5(tensorGemm_io_inp_rd_data_bits_0_5),
    .io_inp_rd_data_bits_0_6(tensorGemm_io_inp_rd_data_bits_0_6),
    .io_inp_rd_data_bits_0_7(tensorGemm_io_inp_rd_data_bits_0_7),
    .io_inp_rd_data_bits_0_8(tensorGemm_io_inp_rd_data_bits_0_8),
    .io_inp_rd_data_bits_0_9(tensorGemm_io_inp_rd_data_bits_0_9),
    .io_inp_rd_data_bits_0_10(tensorGemm_io_inp_rd_data_bits_0_10),
    .io_inp_rd_data_bits_0_11(tensorGemm_io_inp_rd_data_bits_0_11),
    .io_inp_rd_data_bits_0_12(tensorGemm_io_inp_rd_data_bits_0_12),
    .io_inp_rd_data_bits_0_13(tensorGemm_io_inp_rd_data_bits_0_13),
    .io_inp_rd_data_bits_0_14(tensorGemm_io_inp_rd_data_bits_0_14),
    .io_inp_rd_data_bits_0_15(tensorGemm_io_inp_rd_data_bits_0_15),
    .io_wgt_rd_idx_valid(tensorGemm_io_wgt_rd_idx_valid),
    .io_wgt_rd_idx_bits(tensorGemm_io_wgt_rd_idx_bits),
    .io_wgt_rd_data_valid(tensorGemm_io_wgt_rd_data_valid),
    .io_wgt_rd_data_bits_0_0(tensorGemm_io_wgt_rd_data_bits_0_0),
    .io_wgt_rd_data_bits_0_1(tensorGemm_io_wgt_rd_data_bits_0_1),
    .io_wgt_rd_data_bits_0_2(tensorGemm_io_wgt_rd_data_bits_0_2),
    .io_wgt_rd_data_bits_0_3(tensorGemm_io_wgt_rd_data_bits_0_3),
    .io_wgt_rd_data_bits_0_4(tensorGemm_io_wgt_rd_data_bits_0_4),
    .io_wgt_rd_data_bits_0_5(tensorGemm_io_wgt_rd_data_bits_0_5),
    .io_wgt_rd_data_bits_0_6(tensorGemm_io_wgt_rd_data_bits_0_6),
    .io_wgt_rd_data_bits_0_7(tensorGemm_io_wgt_rd_data_bits_0_7),
    .io_wgt_rd_data_bits_0_8(tensorGemm_io_wgt_rd_data_bits_0_8),
    .io_wgt_rd_data_bits_0_9(tensorGemm_io_wgt_rd_data_bits_0_9),
    .io_wgt_rd_data_bits_0_10(tensorGemm_io_wgt_rd_data_bits_0_10),
    .io_wgt_rd_data_bits_0_11(tensorGemm_io_wgt_rd_data_bits_0_11),
    .io_wgt_rd_data_bits_0_12(tensorGemm_io_wgt_rd_data_bits_0_12),
    .io_wgt_rd_data_bits_0_13(tensorGemm_io_wgt_rd_data_bits_0_13),
    .io_wgt_rd_data_bits_0_14(tensorGemm_io_wgt_rd_data_bits_0_14),
    .io_wgt_rd_data_bits_0_15(tensorGemm_io_wgt_rd_data_bits_0_15),
    .io_wgt_rd_data_bits_1_0(tensorGemm_io_wgt_rd_data_bits_1_0),
    .io_wgt_rd_data_bits_1_1(tensorGemm_io_wgt_rd_data_bits_1_1),
    .io_wgt_rd_data_bits_1_2(tensorGemm_io_wgt_rd_data_bits_1_2),
    .io_wgt_rd_data_bits_1_3(tensorGemm_io_wgt_rd_data_bits_1_3),
    .io_wgt_rd_data_bits_1_4(tensorGemm_io_wgt_rd_data_bits_1_4),
    .io_wgt_rd_data_bits_1_5(tensorGemm_io_wgt_rd_data_bits_1_5),
    .io_wgt_rd_data_bits_1_6(tensorGemm_io_wgt_rd_data_bits_1_6),
    .io_wgt_rd_data_bits_1_7(tensorGemm_io_wgt_rd_data_bits_1_7),
    .io_wgt_rd_data_bits_1_8(tensorGemm_io_wgt_rd_data_bits_1_8),
    .io_wgt_rd_data_bits_1_9(tensorGemm_io_wgt_rd_data_bits_1_9),
    .io_wgt_rd_data_bits_1_10(tensorGemm_io_wgt_rd_data_bits_1_10),
    .io_wgt_rd_data_bits_1_11(tensorGemm_io_wgt_rd_data_bits_1_11),
    .io_wgt_rd_data_bits_1_12(tensorGemm_io_wgt_rd_data_bits_1_12),
    .io_wgt_rd_data_bits_1_13(tensorGemm_io_wgt_rd_data_bits_1_13),
    .io_wgt_rd_data_bits_1_14(tensorGemm_io_wgt_rd_data_bits_1_14),
    .io_wgt_rd_data_bits_1_15(tensorGemm_io_wgt_rd_data_bits_1_15),
    .io_wgt_rd_data_bits_2_0(tensorGemm_io_wgt_rd_data_bits_2_0),
    .io_wgt_rd_data_bits_2_1(tensorGemm_io_wgt_rd_data_bits_2_1),
    .io_wgt_rd_data_bits_2_2(tensorGemm_io_wgt_rd_data_bits_2_2),
    .io_wgt_rd_data_bits_2_3(tensorGemm_io_wgt_rd_data_bits_2_3),
    .io_wgt_rd_data_bits_2_4(tensorGemm_io_wgt_rd_data_bits_2_4),
    .io_wgt_rd_data_bits_2_5(tensorGemm_io_wgt_rd_data_bits_2_5),
    .io_wgt_rd_data_bits_2_6(tensorGemm_io_wgt_rd_data_bits_2_6),
    .io_wgt_rd_data_bits_2_7(tensorGemm_io_wgt_rd_data_bits_2_7),
    .io_wgt_rd_data_bits_2_8(tensorGemm_io_wgt_rd_data_bits_2_8),
    .io_wgt_rd_data_bits_2_9(tensorGemm_io_wgt_rd_data_bits_2_9),
    .io_wgt_rd_data_bits_2_10(tensorGemm_io_wgt_rd_data_bits_2_10),
    .io_wgt_rd_data_bits_2_11(tensorGemm_io_wgt_rd_data_bits_2_11),
    .io_wgt_rd_data_bits_2_12(tensorGemm_io_wgt_rd_data_bits_2_12),
    .io_wgt_rd_data_bits_2_13(tensorGemm_io_wgt_rd_data_bits_2_13),
    .io_wgt_rd_data_bits_2_14(tensorGemm_io_wgt_rd_data_bits_2_14),
    .io_wgt_rd_data_bits_2_15(tensorGemm_io_wgt_rd_data_bits_2_15),
    .io_wgt_rd_data_bits_3_0(tensorGemm_io_wgt_rd_data_bits_3_0),
    .io_wgt_rd_data_bits_3_1(tensorGemm_io_wgt_rd_data_bits_3_1),
    .io_wgt_rd_data_bits_3_2(tensorGemm_io_wgt_rd_data_bits_3_2),
    .io_wgt_rd_data_bits_3_3(tensorGemm_io_wgt_rd_data_bits_3_3),
    .io_wgt_rd_data_bits_3_4(tensorGemm_io_wgt_rd_data_bits_3_4),
    .io_wgt_rd_data_bits_3_5(tensorGemm_io_wgt_rd_data_bits_3_5),
    .io_wgt_rd_data_bits_3_6(tensorGemm_io_wgt_rd_data_bits_3_6),
    .io_wgt_rd_data_bits_3_7(tensorGemm_io_wgt_rd_data_bits_3_7),
    .io_wgt_rd_data_bits_3_8(tensorGemm_io_wgt_rd_data_bits_3_8),
    .io_wgt_rd_data_bits_3_9(tensorGemm_io_wgt_rd_data_bits_3_9),
    .io_wgt_rd_data_bits_3_10(tensorGemm_io_wgt_rd_data_bits_3_10),
    .io_wgt_rd_data_bits_3_11(tensorGemm_io_wgt_rd_data_bits_3_11),
    .io_wgt_rd_data_bits_3_12(tensorGemm_io_wgt_rd_data_bits_3_12),
    .io_wgt_rd_data_bits_3_13(tensorGemm_io_wgt_rd_data_bits_3_13),
    .io_wgt_rd_data_bits_3_14(tensorGemm_io_wgt_rd_data_bits_3_14),
    .io_wgt_rd_data_bits_3_15(tensorGemm_io_wgt_rd_data_bits_3_15),
    .io_wgt_rd_data_bits_4_0(tensorGemm_io_wgt_rd_data_bits_4_0),
    .io_wgt_rd_data_bits_4_1(tensorGemm_io_wgt_rd_data_bits_4_1),
    .io_wgt_rd_data_bits_4_2(tensorGemm_io_wgt_rd_data_bits_4_2),
    .io_wgt_rd_data_bits_4_3(tensorGemm_io_wgt_rd_data_bits_4_3),
    .io_wgt_rd_data_bits_4_4(tensorGemm_io_wgt_rd_data_bits_4_4),
    .io_wgt_rd_data_bits_4_5(tensorGemm_io_wgt_rd_data_bits_4_5),
    .io_wgt_rd_data_bits_4_6(tensorGemm_io_wgt_rd_data_bits_4_6),
    .io_wgt_rd_data_bits_4_7(tensorGemm_io_wgt_rd_data_bits_4_7),
    .io_wgt_rd_data_bits_4_8(tensorGemm_io_wgt_rd_data_bits_4_8),
    .io_wgt_rd_data_bits_4_9(tensorGemm_io_wgt_rd_data_bits_4_9),
    .io_wgt_rd_data_bits_4_10(tensorGemm_io_wgt_rd_data_bits_4_10),
    .io_wgt_rd_data_bits_4_11(tensorGemm_io_wgt_rd_data_bits_4_11),
    .io_wgt_rd_data_bits_4_12(tensorGemm_io_wgt_rd_data_bits_4_12),
    .io_wgt_rd_data_bits_4_13(tensorGemm_io_wgt_rd_data_bits_4_13),
    .io_wgt_rd_data_bits_4_14(tensorGemm_io_wgt_rd_data_bits_4_14),
    .io_wgt_rd_data_bits_4_15(tensorGemm_io_wgt_rd_data_bits_4_15),
    .io_wgt_rd_data_bits_5_0(tensorGemm_io_wgt_rd_data_bits_5_0),
    .io_wgt_rd_data_bits_5_1(tensorGemm_io_wgt_rd_data_bits_5_1),
    .io_wgt_rd_data_bits_5_2(tensorGemm_io_wgt_rd_data_bits_5_2),
    .io_wgt_rd_data_bits_5_3(tensorGemm_io_wgt_rd_data_bits_5_3),
    .io_wgt_rd_data_bits_5_4(tensorGemm_io_wgt_rd_data_bits_5_4),
    .io_wgt_rd_data_bits_5_5(tensorGemm_io_wgt_rd_data_bits_5_5),
    .io_wgt_rd_data_bits_5_6(tensorGemm_io_wgt_rd_data_bits_5_6),
    .io_wgt_rd_data_bits_5_7(tensorGemm_io_wgt_rd_data_bits_5_7),
    .io_wgt_rd_data_bits_5_8(tensorGemm_io_wgt_rd_data_bits_5_8),
    .io_wgt_rd_data_bits_5_9(tensorGemm_io_wgt_rd_data_bits_5_9),
    .io_wgt_rd_data_bits_5_10(tensorGemm_io_wgt_rd_data_bits_5_10),
    .io_wgt_rd_data_bits_5_11(tensorGemm_io_wgt_rd_data_bits_5_11),
    .io_wgt_rd_data_bits_5_12(tensorGemm_io_wgt_rd_data_bits_5_12),
    .io_wgt_rd_data_bits_5_13(tensorGemm_io_wgt_rd_data_bits_5_13),
    .io_wgt_rd_data_bits_5_14(tensorGemm_io_wgt_rd_data_bits_5_14),
    .io_wgt_rd_data_bits_5_15(tensorGemm_io_wgt_rd_data_bits_5_15),
    .io_wgt_rd_data_bits_6_0(tensorGemm_io_wgt_rd_data_bits_6_0),
    .io_wgt_rd_data_bits_6_1(tensorGemm_io_wgt_rd_data_bits_6_1),
    .io_wgt_rd_data_bits_6_2(tensorGemm_io_wgt_rd_data_bits_6_2),
    .io_wgt_rd_data_bits_6_3(tensorGemm_io_wgt_rd_data_bits_6_3),
    .io_wgt_rd_data_bits_6_4(tensorGemm_io_wgt_rd_data_bits_6_4),
    .io_wgt_rd_data_bits_6_5(tensorGemm_io_wgt_rd_data_bits_6_5),
    .io_wgt_rd_data_bits_6_6(tensorGemm_io_wgt_rd_data_bits_6_6),
    .io_wgt_rd_data_bits_6_7(tensorGemm_io_wgt_rd_data_bits_6_7),
    .io_wgt_rd_data_bits_6_8(tensorGemm_io_wgt_rd_data_bits_6_8),
    .io_wgt_rd_data_bits_6_9(tensorGemm_io_wgt_rd_data_bits_6_9),
    .io_wgt_rd_data_bits_6_10(tensorGemm_io_wgt_rd_data_bits_6_10),
    .io_wgt_rd_data_bits_6_11(tensorGemm_io_wgt_rd_data_bits_6_11),
    .io_wgt_rd_data_bits_6_12(tensorGemm_io_wgt_rd_data_bits_6_12),
    .io_wgt_rd_data_bits_6_13(tensorGemm_io_wgt_rd_data_bits_6_13),
    .io_wgt_rd_data_bits_6_14(tensorGemm_io_wgt_rd_data_bits_6_14),
    .io_wgt_rd_data_bits_6_15(tensorGemm_io_wgt_rd_data_bits_6_15),
    .io_wgt_rd_data_bits_7_0(tensorGemm_io_wgt_rd_data_bits_7_0),
    .io_wgt_rd_data_bits_7_1(tensorGemm_io_wgt_rd_data_bits_7_1),
    .io_wgt_rd_data_bits_7_2(tensorGemm_io_wgt_rd_data_bits_7_2),
    .io_wgt_rd_data_bits_7_3(tensorGemm_io_wgt_rd_data_bits_7_3),
    .io_wgt_rd_data_bits_7_4(tensorGemm_io_wgt_rd_data_bits_7_4),
    .io_wgt_rd_data_bits_7_5(tensorGemm_io_wgt_rd_data_bits_7_5),
    .io_wgt_rd_data_bits_7_6(tensorGemm_io_wgt_rd_data_bits_7_6),
    .io_wgt_rd_data_bits_7_7(tensorGemm_io_wgt_rd_data_bits_7_7),
    .io_wgt_rd_data_bits_7_8(tensorGemm_io_wgt_rd_data_bits_7_8),
    .io_wgt_rd_data_bits_7_9(tensorGemm_io_wgt_rd_data_bits_7_9),
    .io_wgt_rd_data_bits_7_10(tensorGemm_io_wgt_rd_data_bits_7_10),
    .io_wgt_rd_data_bits_7_11(tensorGemm_io_wgt_rd_data_bits_7_11),
    .io_wgt_rd_data_bits_7_12(tensorGemm_io_wgt_rd_data_bits_7_12),
    .io_wgt_rd_data_bits_7_13(tensorGemm_io_wgt_rd_data_bits_7_13),
    .io_wgt_rd_data_bits_7_14(tensorGemm_io_wgt_rd_data_bits_7_14),
    .io_wgt_rd_data_bits_7_15(tensorGemm_io_wgt_rd_data_bits_7_15),
    .io_wgt_rd_data_bits_8_0(tensorGemm_io_wgt_rd_data_bits_8_0),
    .io_wgt_rd_data_bits_8_1(tensorGemm_io_wgt_rd_data_bits_8_1),
    .io_wgt_rd_data_bits_8_2(tensorGemm_io_wgt_rd_data_bits_8_2),
    .io_wgt_rd_data_bits_8_3(tensorGemm_io_wgt_rd_data_bits_8_3),
    .io_wgt_rd_data_bits_8_4(tensorGemm_io_wgt_rd_data_bits_8_4),
    .io_wgt_rd_data_bits_8_5(tensorGemm_io_wgt_rd_data_bits_8_5),
    .io_wgt_rd_data_bits_8_6(tensorGemm_io_wgt_rd_data_bits_8_6),
    .io_wgt_rd_data_bits_8_7(tensorGemm_io_wgt_rd_data_bits_8_7),
    .io_wgt_rd_data_bits_8_8(tensorGemm_io_wgt_rd_data_bits_8_8),
    .io_wgt_rd_data_bits_8_9(tensorGemm_io_wgt_rd_data_bits_8_9),
    .io_wgt_rd_data_bits_8_10(tensorGemm_io_wgt_rd_data_bits_8_10),
    .io_wgt_rd_data_bits_8_11(tensorGemm_io_wgt_rd_data_bits_8_11),
    .io_wgt_rd_data_bits_8_12(tensorGemm_io_wgt_rd_data_bits_8_12),
    .io_wgt_rd_data_bits_8_13(tensorGemm_io_wgt_rd_data_bits_8_13),
    .io_wgt_rd_data_bits_8_14(tensorGemm_io_wgt_rd_data_bits_8_14),
    .io_wgt_rd_data_bits_8_15(tensorGemm_io_wgt_rd_data_bits_8_15),
    .io_wgt_rd_data_bits_9_0(tensorGemm_io_wgt_rd_data_bits_9_0),
    .io_wgt_rd_data_bits_9_1(tensorGemm_io_wgt_rd_data_bits_9_1),
    .io_wgt_rd_data_bits_9_2(tensorGemm_io_wgt_rd_data_bits_9_2),
    .io_wgt_rd_data_bits_9_3(tensorGemm_io_wgt_rd_data_bits_9_3),
    .io_wgt_rd_data_bits_9_4(tensorGemm_io_wgt_rd_data_bits_9_4),
    .io_wgt_rd_data_bits_9_5(tensorGemm_io_wgt_rd_data_bits_9_5),
    .io_wgt_rd_data_bits_9_6(tensorGemm_io_wgt_rd_data_bits_9_6),
    .io_wgt_rd_data_bits_9_7(tensorGemm_io_wgt_rd_data_bits_9_7),
    .io_wgt_rd_data_bits_9_8(tensorGemm_io_wgt_rd_data_bits_9_8),
    .io_wgt_rd_data_bits_9_9(tensorGemm_io_wgt_rd_data_bits_9_9),
    .io_wgt_rd_data_bits_9_10(tensorGemm_io_wgt_rd_data_bits_9_10),
    .io_wgt_rd_data_bits_9_11(tensorGemm_io_wgt_rd_data_bits_9_11),
    .io_wgt_rd_data_bits_9_12(tensorGemm_io_wgt_rd_data_bits_9_12),
    .io_wgt_rd_data_bits_9_13(tensorGemm_io_wgt_rd_data_bits_9_13),
    .io_wgt_rd_data_bits_9_14(tensorGemm_io_wgt_rd_data_bits_9_14),
    .io_wgt_rd_data_bits_9_15(tensorGemm_io_wgt_rd_data_bits_9_15),
    .io_wgt_rd_data_bits_10_0(tensorGemm_io_wgt_rd_data_bits_10_0),
    .io_wgt_rd_data_bits_10_1(tensorGemm_io_wgt_rd_data_bits_10_1),
    .io_wgt_rd_data_bits_10_2(tensorGemm_io_wgt_rd_data_bits_10_2),
    .io_wgt_rd_data_bits_10_3(tensorGemm_io_wgt_rd_data_bits_10_3),
    .io_wgt_rd_data_bits_10_4(tensorGemm_io_wgt_rd_data_bits_10_4),
    .io_wgt_rd_data_bits_10_5(tensorGemm_io_wgt_rd_data_bits_10_5),
    .io_wgt_rd_data_bits_10_6(tensorGemm_io_wgt_rd_data_bits_10_6),
    .io_wgt_rd_data_bits_10_7(tensorGemm_io_wgt_rd_data_bits_10_7),
    .io_wgt_rd_data_bits_10_8(tensorGemm_io_wgt_rd_data_bits_10_8),
    .io_wgt_rd_data_bits_10_9(tensorGemm_io_wgt_rd_data_bits_10_9),
    .io_wgt_rd_data_bits_10_10(tensorGemm_io_wgt_rd_data_bits_10_10),
    .io_wgt_rd_data_bits_10_11(tensorGemm_io_wgt_rd_data_bits_10_11),
    .io_wgt_rd_data_bits_10_12(tensorGemm_io_wgt_rd_data_bits_10_12),
    .io_wgt_rd_data_bits_10_13(tensorGemm_io_wgt_rd_data_bits_10_13),
    .io_wgt_rd_data_bits_10_14(tensorGemm_io_wgt_rd_data_bits_10_14),
    .io_wgt_rd_data_bits_10_15(tensorGemm_io_wgt_rd_data_bits_10_15),
    .io_wgt_rd_data_bits_11_0(tensorGemm_io_wgt_rd_data_bits_11_0),
    .io_wgt_rd_data_bits_11_1(tensorGemm_io_wgt_rd_data_bits_11_1),
    .io_wgt_rd_data_bits_11_2(tensorGemm_io_wgt_rd_data_bits_11_2),
    .io_wgt_rd_data_bits_11_3(tensorGemm_io_wgt_rd_data_bits_11_3),
    .io_wgt_rd_data_bits_11_4(tensorGemm_io_wgt_rd_data_bits_11_4),
    .io_wgt_rd_data_bits_11_5(tensorGemm_io_wgt_rd_data_bits_11_5),
    .io_wgt_rd_data_bits_11_6(tensorGemm_io_wgt_rd_data_bits_11_6),
    .io_wgt_rd_data_bits_11_7(tensorGemm_io_wgt_rd_data_bits_11_7),
    .io_wgt_rd_data_bits_11_8(tensorGemm_io_wgt_rd_data_bits_11_8),
    .io_wgt_rd_data_bits_11_9(tensorGemm_io_wgt_rd_data_bits_11_9),
    .io_wgt_rd_data_bits_11_10(tensorGemm_io_wgt_rd_data_bits_11_10),
    .io_wgt_rd_data_bits_11_11(tensorGemm_io_wgt_rd_data_bits_11_11),
    .io_wgt_rd_data_bits_11_12(tensorGemm_io_wgt_rd_data_bits_11_12),
    .io_wgt_rd_data_bits_11_13(tensorGemm_io_wgt_rd_data_bits_11_13),
    .io_wgt_rd_data_bits_11_14(tensorGemm_io_wgt_rd_data_bits_11_14),
    .io_wgt_rd_data_bits_11_15(tensorGemm_io_wgt_rd_data_bits_11_15),
    .io_wgt_rd_data_bits_12_0(tensorGemm_io_wgt_rd_data_bits_12_0),
    .io_wgt_rd_data_bits_12_1(tensorGemm_io_wgt_rd_data_bits_12_1),
    .io_wgt_rd_data_bits_12_2(tensorGemm_io_wgt_rd_data_bits_12_2),
    .io_wgt_rd_data_bits_12_3(tensorGemm_io_wgt_rd_data_bits_12_3),
    .io_wgt_rd_data_bits_12_4(tensorGemm_io_wgt_rd_data_bits_12_4),
    .io_wgt_rd_data_bits_12_5(tensorGemm_io_wgt_rd_data_bits_12_5),
    .io_wgt_rd_data_bits_12_6(tensorGemm_io_wgt_rd_data_bits_12_6),
    .io_wgt_rd_data_bits_12_7(tensorGemm_io_wgt_rd_data_bits_12_7),
    .io_wgt_rd_data_bits_12_8(tensorGemm_io_wgt_rd_data_bits_12_8),
    .io_wgt_rd_data_bits_12_9(tensorGemm_io_wgt_rd_data_bits_12_9),
    .io_wgt_rd_data_bits_12_10(tensorGemm_io_wgt_rd_data_bits_12_10),
    .io_wgt_rd_data_bits_12_11(tensorGemm_io_wgt_rd_data_bits_12_11),
    .io_wgt_rd_data_bits_12_12(tensorGemm_io_wgt_rd_data_bits_12_12),
    .io_wgt_rd_data_bits_12_13(tensorGemm_io_wgt_rd_data_bits_12_13),
    .io_wgt_rd_data_bits_12_14(tensorGemm_io_wgt_rd_data_bits_12_14),
    .io_wgt_rd_data_bits_12_15(tensorGemm_io_wgt_rd_data_bits_12_15),
    .io_wgt_rd_data_bits_13_0(tensorGemm_io_wgt_rd_data_bits_13_0),
    .io_wgt_rd_data_bits_13_1(tensorGemm_io_wgt_rd_data_bits_13_1),
    .io_wgt_rd_data_bits_13_2(tensorGemm_io_wgt_rd_data_bits_13_2),
    .io_wgt_rd_data_bits_13_3(tensorGemm_io_wgt_rd_data_bits_13_3),
    .io_wgt_rd_data_bits_13_4(tensorGemm_io_wgt_rd_data_bits_13_4),
    .io_wgt_rd_data_bits_13_5(tensorGemm_io_wgt_rd_data_bits_13_5),
    .io_wgt_rd_data_bits_13_6(tensorGemm_io_wgt_rd_data_bits_13_6),
    .io_wgt_rd_data_bits_13_7(tensorGemm_io_wgt_rd_data_bits_13_7),
    .io_wgt_rd_data_bits_13_8(tensorGemm_io_wgt_rd_data_bits_13_8),
    .io_wgt_rd_data_bits_13_9(tensorGemm_io_wgt_rd_data_bits_13_9),
    .io_wgt_rd_data_bits_13_10(tensorGemm_io_wgt_rd_data_bits_13_10),
    .io_wgt_rd_data_bits_13_11(tensorGemm_io_wgt_rd_data_bits_13_11),
    .io_wgt_rd_data_bits_13_12(tensorGemm_io_wgt_rd_data_bits_13_12),
    .io_wgt_rd_data_bits_13_13(tensorGemm_io_wgt_rd_data_bits_13_13),
    .io_wgt_rd_data_bits_13_14(tensorGemm_io_wgt_rd_data_bits_13_14),
    .io_wgt_rd_data_bits_13_15(tensorGemm_io_wgt_rd_data_bits_13_15),
    .io_wgt_rd_data_bits_14_0(tensorGemm_io_wgt_rd_data_bits_14_0),
    .io_wgt_rd_data_bits_14_1(tensorGemm_io_wgt_rd_data_bits_14_1),
    .io_wgt_rd_data_bits_14_2(tensorGemm_io_wgt_rd_data_bits_14_2),
    .io_wgt_rd_data_bits_14_3(tensorGemm_io_wgt_rd_data_bits_14_3),
    .io_wgt_rd_data_bits_14_4(tensorGemm_io_wgt_rd_data_bits_14_4),
    .io_wgt_rd_data_bits_14_5(tensorGemm_io_wgt_rd_data_bits_14_5),
    .io_wgt_rd_data_bits_14_6(tensorGemm_io_wgt_rd_data_bits_14_6),
    .io_wgt_rd_data_bits_14_7(tensorGemm_io_wgt_rd_data_bits_14_7),
    .io_wgt_rd_data_bits_14_8(tensorGemm_io_wgt_rd_data_bits_14_8),
    .io_wgt_rd_data_bits_14_9(tensorGemm_io_wgt_rd_data_bits_14_9),
    .io_wgt_rd_data_bits_14_10(tensorGemm_io_wgt_rd_data_bits_14_10),
    .io_wgt_rd_data_bits_14_11(tensorGemm_io_wgt_rd_data_bits_14_11),
    .io_wgt_rd_data_bits_14_12(tensorGemm_io_wgt_rd_data_bits_14_12),
    .io_wgt_rd_data_bits_14_13(tensorGemm_io_wgt_rd_data_bits_14_13),
    .io_wgt_rd_data_bits_14_14(tensorGemm_io_wgt_rd_data_bits_14_14),
    .io_wgt_rd_data_bits_14_15(tensorGemm_io_wgt_rd_data_bits_14_15),
    .io_wgt_rd_data_bits_15_0(tensorGemm_io_wgt_rd_data_bits_15_0),
    .io_wgt_rd_data_bits_15_1(tensorGemm_io_wgt_rd_data_bits_15_1),
    .io_wgt_rd_data_bits_15_2(tensorGemm_io_wgt_rd_data_bits_15_2),
    .io_wgt_rd_data_bits_15_3(tensorGemm_io_wgt_rd_data_bits_15_3),
    .io_wgt_rd_data_bits_15_4(tensorGemm_io_wgt_rd_data_bits_15_4),
    .io_wgt_rd_data_bits_15_5(tensorGemm_io_wgt_rd_data_bits_15_5),
    .io_wgt_rd_data_bits_15_6(tensorGemm_io_wgt_rd_data_bits_15_6),
    .io_wgt_rd_data_bits_15_7(tensorGemm_io_wgt_rd_data_bits_15_7),
    .io_wgt_rd_data_bits_15_8(tensorGemm_io_wgt_rd_data_bits_15_8),
    .io_wgt_rd_data_bits_15_9(tensorGemm_io_wgt_rd_data_bits_15_9),
    .io_wgt_rd_data_bits_15_10(tensorGemm_io_wgt_rd_data_bits_15_10),
    .io_wgt_rd_data_bits_15_11(tensorGemm_io_wgt_rd_data_bits_15_11),
    .io_wgt_rd_data_bits_15_12(tensorGemm_io_wgt_rd_data_bits_15_12),
    .io_wgt_rd_data_bits_15_13(tensorGemm_io_wgt_rd_data_bits_15_13),
    .io_wgt_rd_data_bits_15_14(tensorGemm_io_wgt_rd_data_bits_15_14),
    .io_wgt_rd_data_bits_15_15(tensorGemm_io_wgt_rd_data_bits_15_15),
    .io_acc_rd_idx_valid(tensorGemm_io_acc_rd_idx_valid),
    .io_acc_rd_idx_bits(tensorGemm_io_acc_rd_idx_bits),
    .io_acc_rd_data_valid(tensorGemm_io_acc_rd_data_valid),
    .io_acc_rd_data_bits_0_0(tensorGemm_io_acc_rd_data_bits_0_0),
    .io_acc_rd_data_bits_0_1(tensorGemm_io_acc_rd_data_bits_0_1),
    .io_acc_rd_data_bits_0_2(tensorGemm_io_acc_rd_data_bits_0_2),
    .io_acc_rd_data_bits_0_3(tensorGemm_io_acc_rd_data_bits_0_3),
    .io_acc_rd_data_bits_0_4(tensorGemm_io_acc_rd_data_bits_0_4),
    .io_acc_rd_data_bits_0_5(tensorGemm_io_acc_rd_data_bits_0_5),
    .io_acc_rd_data_bits_0_6(tensorGemm_io_acc_rd_data_bits_0_6),
    .io_acc_rd_data_bits_0_7(tensorGemm_io_acc_rd_data_bits_0_7),
    .io_acc_rd_data_bits_0_8(tensorGemm_io_acc_rd_data_bits_0_8),
    .io_acc_rd_data_bits_0_9(tensorGemm_io_acc_rd_data_bits_0_9),
    .io_acc_rd_data_bits_0_10(tensorGemm_io_acc_rd_data_bits_0_10),
    .io_acc_rd_data_bits_0_11(tensorGemm_io_acc_rd_data_bits_0_11),
    .io_acc_rd_data_bits_0_12(tensorGemm_io_acc_rd_data_bits_0_12),
    .io_acc_rd_data_bits_0_13(tensorGemm_io_acc_rd_data_bits_0_13),
    .io_acc_rd_data_bits_0_14(tensorGemm_io_acc_rd_data_bits_0_14),
    .io_acc_rd_data_bits_0_15(tensorGemm_io_acc_rd_data_bits_0_15),
    .io_acc_wr_valid(tensorGemm_io_acc_wr_valid),
    .io_acc_wr_bits_idx(tensorGemm_io_acc_wr_bits_idx),
    .io_acc_wr_bits_data_0_0(tensorGemm_io_acc_wr_bits_data_0_0),
    .io_acc_wr_bits_data_0_1(tensorGemm_io_acc_wr_bits_data_0_1),
    .io_acc_wr_bits_data_0_2(tensorGemm_io_acc_wr_bits_data_0_2),
    .io_acc_wr_bits_data_0_3(tensorGemm_io_acc_wr_bits_data_0_3),
    .io_acc_wr_bits_data_0_4(tensorGemm_io_acc_wr_bits_data_0_4),
    .io_acc_wr_bits_data_0_5(tensorGemm_io_acc_wr_bits_data_0_5),
    .io_acc_wr_bits_data_0_6(tensorGemm_io_acc_wr_bits_data_0_6),
    .io_acc_wr_bits_data_0_7(tensorGemm_io_acc_wr_bits_data_0_7),
    .io_acc_wr_bits_data_0_8(tensorGemm_io_acc_wr_bits_data_0_8),
    .io_acc_wr_bits_data_0_9(tensorGemm_io_acc_wr_bits_data_0_9),
    .io_acc_wr_bits_data_0_10(tensorGemm_io_acc_wr_bits_data_0_10),
    .io_acc_wr_bits_data_0_11(tensorGemm_io_acc_wr_bits_data_0_11),
    .io_acc_wr_bits_data_0_12(tensorGemm_io_acc_wr_bits_data_0_12),
    .io_acc_wr_bits_data_0_13(tensorGemm_io_acc_wr_bits_data_0_13),
    .io_acc_wr_bits_data_0_14(tensorGemm_io_acc_wr_bits_data_0_14),
    .io_acc_wr_bits_data_0_15(tensorGemm_io_acc_wr_bits_data_0_15),
    .io_out_wr_valid(tensorGemm_io_out_wr_valid),
    .io_out_wr_bits_idx(tensorGemm_io_out_wr_bits_idx),
    .io_out_wr_bits_data_0_0(tensorGemm_io_out_wr_bits_data_0_0),
    .io_out_wr_bits_data_0_1(tensorGemm_io_out_wr_bits_data_0_1),
    .io_out_wr_bits_data_0_2(tensorGemm_io_out_wr_bits_data_0_2),
    .io_out_wr_bits_data_0_3(tensorGemm_io_out_wr_bits_data_0_3),
    .io_out_wr_bits_data_0_4(tensorGemm_io_out_wr_bits_data_0_4),
    .io_out_wr_bits_data_0_5(tensorGemm_io_out_wr_bits_data_0_5),
    .io_out_wr_bits_data_0_6(tensorGemm_io_out_wr_bits_data_0_6),
    .io_out_wr_bits_data_0_7(tensorGemm_io_out_wr_bits_data_0_7),
    .io_out_wr_bits_data_0_8(tensorGemm_io_out_wr_bits_data_0_8),
    .io_out_wr_bits_data_0_9(tensorGemm_io_out_wr_bits_data_0_9),
    .io_out_wr_bits_data_0_10(tensorGemm_io_out_wr_bits_data_0_10),
    .io_out_wr_bits_data_0_11(tensorGemm_io_out_wr_bits_data_0_11),
    .io_out_wr_bits_data_0_12(tensorGemm_io_out_wr_bits_data_0_12),
    .io_out_wr_bits_data_0_13(tensorGemm_io_out_wr_bits_data_0_13),
    .io_out_wr_bits_data_0_14(tensorGemm_io_out_wr_bits_data_0_14),
    .io_out_wr_bits_data_0_15(tensorGemm_io_out_wr_bits_data_0_15)
  );
  TensorAlu tensorAlu ( // @[Compute.scala 59:25:@23209.4]
    .clock(tensorAlu_clock),
    .reset(tensorAlu_reset),
    .io_start(tensorAlu_io_start),
    .io_done(tensorAlu_io_done),
    .io_inst(tensorAlu_io_inst),
    .io_uop_idx_valid(tensorAlu_io_uop_idx_valid),
    .io_uop_idx_bits(tensorAlu_io_uop_idx_bits),
    .io_uop_data_valid(tensorAlu_io_uop_data_valid),
    .io_uop_data_bits_u1(tensorAlu_io_uop_data_bits_u1),
    .io_uop_data_bits_u0(tensorAlu_io_uop_data_bits_u0),
    .io_acc_rd_idx_valid(tensorAlu_io_acc_rd_idx_valid),
    .io_acc_rd_idx_bits(tensorAlu_io_acc_rd_idx_bits),
    .io_acc_rd_data_valid(tensorAlu_io_acc_rd_data_valid),
    .io_acc_rd_data_bits_0_0(tensorAlu_io_acc_rd_data_bits_0_0),
    .io_acc_rd_data_bits_0_1(tensorAlu_io_acc_rd_data_bits_0_1),
    .io_acc_rd_data_bits_0_2(tensorAlu_io_acc_rd_data_bits_0_2),
    .io_acc_rd_data_bits_0_3(tensorAlu_io_acc_rd_data_bits_0_3),
    .io_acc_rd_data_bits_0_4(tensorAlu_io_acc_rd_data_bits_0_4),
    .io_acc_rd_data_bits_0_5(tensorAlu_io_acc_rd_data_bits_0_5),
    .io_acc_rd_data_bits_0_6(tensorAlu_io_acc_rd_data_bits_0_6),
    .io_acc_rd_data_bits_0_7(tensorAlu_io_acc_rd_data_bits_0_7),
    .io_acc_rd_data_bits_0_8(tensorAlu_io_acc_rd_data_bits_0_8),
    .io_acc_rd_data_bits_0_9(tensorAlu_io_acc_rd_data_bits_0_9),
    .io_acc_rd_data_bits_0_10(tensorAlu_io_acc_rd_data_bits_0_10),
    .io_acc_rd_data_bits_0_11(tensorAlu_io_acc_rd_data_bits_0_11),
    .io_acc_rd_data_bits_0_12(tensorAlu_io_acc_rd_data_bits_0_12),
    .io_acc_rd_data_bits_0_13(tensorAlu_io_acc_rd_data_bits_0_13),
    .io_acc_rd_data_bits_0_14(tensorAlu_io_acc_rd_data_bits_0_14),
    .io_acc_rd_data_bits_0_15(tensorAlu_io_acc_rd_data_bits_0_15),
    .io_acc_wr_valid(tensorAlu_io_acc_wr_valid),
    .io_acc_wr_bits_idx(tensorAlu_io_acc_wr_bits_idx),
    .io_acc_wr_bits_data_0_0(tensorAlu_io_acc_wr_bits_data_0_0),
    .io_acc_wr_bits_data_0_1(tensorAlu_io_acc_wr_bits_data_0_1),
    .io_acc_wr_bits_data_0_2(tensorAlu_io_acc_wr_bits_data_0_2),
    .io_acc_wr_bits_data_0_3(tensorAlu_io_acc_wr_bits_data_0_3),
    .io_acc_wr_bits_data_0_4(tensorAlu_io_acc_wr_bits_data_0_4),
    .io_acc_wr_bits_data_0_5(tensorAlu_io_acc_wr_bits_data_0_5),
    .io_acc_wr_bits_data_0_6(tensorAlu_io_acc_wr_bits_data_0_6),
    .io_acc_wr_bits_data_0_7(tensorAlu_io_acc_wr_bits_data_0_7),
    .io_acc_wr_bits_data_0_8(tensorAlu_io_acc_wr_bits_data_0_8),
    .io_acc_wr_bits_data_0_9(tensorAlu_io_acc_wr_bits_data_0_9),
    .io_acc_wr_bits_data_0_10(tensorAlu_io_acc_wr_bits_data_0_10),
    .io_acc_wr_bits_data_0_11(tensorAlu_io_acc_wr_bits_data_0_11),
    .io_acc_wr_bits_data_0_12(tensorAlu_io_acc_wr_bits_data_0_12),
    .io_acc_wr_bits_data_0_13(tensorAlu_io_acc_wr_bits_data_0_13),
    .io_acc_wr_bits_data_0_14(tensorAlu_io_acc_wr_bits_data_0_14),
    .io_acc_wr_bits_data_0_15(tensorAlu_io_acc_wr_bits_data_0_15),
    .io_out_wr_valid(tensorAlu_io_out_wr_valid),
    .io_out_wr_bits_idx(tensorAlu_io_out_wr_bits_idx),
    .io_out_wr_bits_data_0_0(tensorAlu_io_out_wr_bits_data_0_0),
    .io_out_wr_bits_data_0_1(tensorAlu_io_out_wr_bits_data_0_1),
    .io_out_wr_bits_data_0_2(tensorAlu_io_out_wr_bits_data_0_2),
    .io_out_wr_bits_data_0_3(tensorAlu_io_out_wr_bits_data_0_3),
    .io_out_wr_bits_data_0_4(tensorAlu_io_out_wr_bits_data_0_4),
    .io_out_wr_bits_data_0_5(tensorAlu_io_out_wr_bits_data_0_5),
    .io_out_wr_bits_data_0_6(tensorAlu_io_out_wr_bits_data_0_6),
    .io_out_wr_bits_data_0_7(tensorAlu_io_out_wr_bits_data_0_7),
    .io_out_wr_bits_data_0_8(tensorAlu_io_out_wr_bits_data_0_8),
    .io_out_wr_bits_data_0_9(tensorAlu_io_out_wr_bits_data_0_9),
    .io_out_wr_bits_data_0_10(tensorAlu_io_out_wr_bits_data_0_10),
    .io_out_wr_bits_data_0_11(tensorAlu_io_out_wr_bits_data_0_11),
    .io_out_wr_bits_data_0_12(tensorAlu_io_out_wr_bits_data_0_12),
    .io_out_wr_bits_data_0_13(tensorAlu_io_out_wr_bits_data_0_13),
    .io_out_wr_bits_data_0_14(tensorAlu_io_out_wr_bits_data_0_14),
    .io_out_wr_bits_data_0_15(tensorAlu_io_out_wr_bits_data_0_15)
  );
  Queue_1 inst_q ( // @[Compute.scala 61:22:@23212.4]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits)
  );
  ComputeDecode dec ( // @[Compute.scala 64:19:@23215.4]
    .io_inst(dec_io_inst),
    .io_push_next(dec_io_push_next),
    .io_push_prev(dec_io_push_prev),
    .io_pop_next(dec_io_pop_next),
    .io_pop_prev(dec_io_pop_prev),
    .io_isLoadAcc(dec_io_isLoadAcc),
    .io_isLoadUop(dec_io_isLoadUop),
    .io_isSync(dec_io_isSync),
    .io_isAlu(dec_io_isAlu),
    .io_isGemm(dec_io_isGemm),
    .io_isFinish(dec_io_isFinish)
  );
  assign inst_type = {dec_io_isFinish,dec_io_isAlu,dec_io_isGemm,dec_io_isLoadAcc,dec_io_isLoadUop}; // @[Cat.scala 30:58:@23222.4]
  assign _T_7054 = dec_io_pop_prev ? s_0_io_sready : 1'h1; // @[Compute.scala 74:40:@23223.4]
  assign sprev = inst_q_io_deq_valid & _T_7054; // @[Compute.scala 74:35:@23224.4]
  assign _T_7056 = dec_io_pop_next ? s_1_io_sready : 1'h1; // @[Compute.scala 75:40:@23225.4]
  assign snext = inst_q_io_deq_valid & _T_7056; // @[Compute.scala 75:35:@23226.4]
  assign start = snext & sprev; // @[Compute.scala 76:21:@23227.4]
  assign _T_7064 = 5'h10 == inst_type; // @[Mux.scala 46:19:@23228.4]
  assign _T_7066 = 5'h8 == inst_type; // @[Mux.scala 46:19:@23230.4]
  assign _T_7067 = _T_7066 ? tensorAlu_io_done : _T_7064; // @[Mux.scala 46:16:@23231.4]
  assign _T_7068 = 5'h4 == inst_type; // @[Mux.scala 46:19:@23232.4]
  assign _T_7069 = _T_7068 ? tensorGemm_io_done : _T_7067; // @[Mux.scala 46:16:@23233.4]
  assign _T_7070 = 5'h2 == inst_type; // @[Mux.scala 46:19:@23234.4]
  assign _T_7071 = _T_7070 ? tensorAcc_io_done : _T_7069; // @[Mux.scala 46:16:@23235.4]
  assign _T_7072 = 5'h1 == inst_type; // @[Mux.scala 46:19:@23236.4]
  assign done = _T_7072 ? loadUop_io_done : _T_7071; // @[Mux.scala 46:16:@23237.4]
  assign _T_7073 = 2'h0 == state; // @[Conditional.scala 37:30:@23238.4]
  assign _T_7075 = inst_type != 5'h0; // @[Compute.scala 96:30:@23245.10]
  assign _GEN_0 = _T_7075 ? 2'h2 : state; // @[Compute.scala 96:35:@23246.10]
  assign _GEN_1 = dec_io_isSync ? 2'h1 : _GEN_0; // @[Compute.scala 94:29:@23241.8]
  assign _GEN_2 = start ? _GEN_1 : state; // @[Compute.scala 93:19:@23240.6]
  assign _T_7076 = 2'h1 == state; // @[Conditional.scala 37:30:@23252.6]
  assign _T_7077 = 2'h2 == state; // @[Conditional.scala 37:30:@23257.8]
  assign _GEN_3 = done ? 2'h0 : state; // @[Compute.scala 105:18:@23259.10]
  assign _GEN_4 = _T_7077 ? _GEN_3 : state; // @[Conditional.scala 39:67:@23258.8]
  assign _GEN_5 = _T_7076 ? 2'h0 : _GEN_4; // @[Conditional.scala 39:67:@23253.6]
  assign _GEN_6 = _T_7073 ? _GEN_2 : _GEN_5; // @[Conditional.scala 40:58:@23239.4]
  assign _T_7078 = state == 2'h2; // @[Compute.scala 113:33:@23266.4]
  assign _T_7079 = _T_7078 & done; // @[Compute.scala 113:42:@23267.4]
  assign _T_7080 = state == 2'h1; // @[Compute.scala 113:59:@23268.4]
  assign _T_7081 = _T_7079 | _T_7080; // @[Compute.scala 113:50:@23269.4]
  assign _T_7082 = state == 2'h0; // @[Compute.scala 116:29:@23271.4]
  assign _T_7083 = _T_7082 & start; // @[Compute.scala 116:39:@23272.4]
  assign io_o_post_0 = dec_io_push_prev & _T_7081; // @[Compute.scala 164:16:@24006.4]
  assign io_o_post_1 = dec_io_push_next & _T_7081; // @[Compute.scala 165:16:@24012.4]
  assign io_inst_ready = inst_q_io_enq_ready; // @[Compute.scala 112:17:@23265.4]
  assign io_vme_rd_0_cmd_valid = loadUop_io_vme_rd_cmd_valid; // @[Compute.scala 119:16:@23282.4]
  assign io_vme_rd_0_cmd_bits_addr = loadUop_io_vme_rd_cmd_bits_addr; // @[Compute.scala 119:16:@23281.4]
  assign io_vme_rd_0_cmd_bits_len = loadUop_io_vme_rd_cmd_bits_len; // @[Compute.scala 119:16:@23280.4]
  assign io_vme_rd_0_data_ready = loadUop_io_vme_rd_data_ready; // @[Compute.scala 119:16:@23279.4]
  assign io_vme_rd_1_cmd_valid = tensorAcc_io_vme_rd_cmd_valid; // @[Compute.scala 128:16:@23320.4]
  assign io_vme_rd_1_cmd_bits_addr = tensorAcc_io_vme_rd_cmd_bits_addr; // @[Compute.scala 128:16:@23319.4]
  assign io_vme_rd_1_cmd_bits_len = tensorAcc_io_vme_rd_cmd_bits_len; // @[Compute.scala 128:16:@23318.4]
  assign io_vme_rd_1_data_ready = tensorAcc_io_vme_rd_data_ready; // @[Compute.scala 128:16:@23317.4]
  assign io_inp_rd_idx_valid = tensorGemm_io_inp_rd_idx_valid; // @[Compute.scala 136:21:@23369.4]
  assign io_inp_rd_idx_bits = tensorGemm_io_inp_rd_idx_bits; // @[Compute.scala 136:21:@23368.4]
  assign io_wgt_rd_idx_valid = tensorGemm_io_wgt_rd_idx_valid; // @[Compute.scala 137:21:@23886.4]
  assign io_wgt_rd_idx_bits = tensorGemm_io_wgt_rd_idx_bits; // @[Compute.scala 137:21:@23885.4]
  assign io_out_wr_valid = dec_io_isGemm ? tensorGemm_io_out_wr_valid : tensorAlu_io_out_wr_valid; // @[Compute.scala 157:13:@23990.4]
  assign io_out_wr_bits_idx = dec_io_isGemm ? tensorGemm_io_out_wr_bits_idx : tensorAlu_io_out_wr_bits_idx; // @[Compute.scala 157:13:@23989.4]
  assign io_out_wr_bits_data_0_0 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_0 : tensorAlu_io_out_wr_bits_data_0_0; // @[Compute.scala 157:13:@23973.4]
  assign io_out_wr_bits_data_0_1 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_1 : tensorAlu_io_out_wr_bits_data_0_1; // @[Compute.scala 157:13:@23974.4]
  assign io_out_wr_bits_data_0_2 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_2 : tensorAlu_io_out_wr_bits_data_0_2; // @[Compute.scala 157:13:@23975.4]
  assign io_out_wr_bits_data_0_3 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_3 : tensorAlu_io_out_wr_bits_data_0_3; // @[Compute.scala 157:13:@23976.4]
  assign io_out_wr_bits_data_0_4 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_4 : tensorAlu_io_out_wr_bits_data_0_4; // @[Compute.scala 157:13:@23977.4]
  assign io_out_wr_bits_data_0_5 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_5 : tensorAlu_io_out_wr_bits_data_0_5; // @[Compute.scala 157:13:@23978.4]
  assign io_out_wr_bits_data_0_6 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_6 : tensorAlu_io_out_wr_bits_data_0_6; // @[Compute.scala 157:13:@23979.4]
  assign io_out_wr_bits_data_0_7 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_7 : tensorAlu_io_out_wr_bits_data_0_7; // @[Compute.scala 157:13:@23980.4]
  assign io_out_wr_bits_data_0_8 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_8 : tensorAlu_io_out_wr_bits_data_0_8; // @[Compute.scala 157:13:@23981.4]
  assign io_out_wr_bits_data_0_9 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_9 : tensorAlu_io_out_wr_bits_data_0_9; // @[Compute.scala 157:13:@23982.4]
  assign io_out_wr_bits_data_0_10 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_10 : tensorAlu_io_out_wr_bits_data_0_10; // @[Compute.scala 157:13:@23983.4]
  assign io_out_wr_bits_data_0_11 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_11 : tensorAlu_io_out_wr_bits_data_0_11; // @[Compute.scala 157:13:@23984.4]
  assign io_out_wr_bits_data_0_12 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_12 : tensorAlu_io_out_wr_bits_data_0_12; // @[Compute.scala 157:13:@23985.4]
  assign io_out_wr_bits_data_0_13 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_13 : tensorAlu_io_out_wr_bits_data_0_13; // @[Compute.scala 157:13:@23986.4]
  assign io_out_wr_bits_data_0_14 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_14 : tensorAlu_io_out_wr_bits_data_0_14; // @[Compute.scala 157:13:@23987.4]
  assign io_out_wr_bits_data_0_15 = dec_io_isGemm ? tensorGemm_io_out_wr_bits_data_0_15 : tensorAlu_io_out_wr_bits_data_0_15; // @[Compute.scala 157:13:@23988.4]
  assign io_finish = _T_7079 & dec_io_isFinish; // @[Compute.scala 168:13:@24016.4]
  assign io_acc_wr_event = tensorAcc_io_tensor_wr_valid; // @[Compute.scala 129:19:@23322.4]
  assign s_0_clock = clock; // @[:@23195.4]
  assign s_0_reset = reset; // @[:@23196.4]
  assign s_0_io_spost = io_i_post_0; // @[Compute.scala 160:17:@23991.4]
  assign s_0_io_swait = dec_io_pop_prev & _T_7083; // @[Compute.scala 162:17:@23996.4]
  assign s_1_clock = clock; // @[:@23198.4]
  assign s_1_reset = reset; // @[:@23199.4]
  assign s_1_io_spost = io_i_post_1; // @[Compute.scala 161:17:@23992.4]
  assign s_1_io_swait = dec_io_pop_next & _T_7083; // @[Compute.scala 163:17:@24000.4]
  assign loadUop_clock = clock; // @[:@23201.4]
  assign loadUop_reset = reset; // @[:@23202.4]
  assign loadUop_io_start = _T_7083 & dec_io_isLoadUop; // @[Compute.scala 116:20:@23274.4]
  assign loadUop_io_inst = inst_q_io_deq_bits; // @[Compute.scala 117:19:@23275.4]
  assign loadUop_io_baddr = io_uop_baddr; // @[Compute.scala 118:20:@23276.4]
  assign loadUop_io_vme_rd_cmd_ready = io_vme_rd_0_cmd_ready; // @[Compute.scala 119:16:@23283.4]
  assign loadUop_io_vme_rd_data_valid = io_vme_rd_0_data_valid; // @[Compute.scala 119:16:@23278.4]
  assign loadUop_io_vme_rd_data_bits = io_vme_rd_0_data_bits; // @[Compute.scala 119:16:@23277.4]
  assign loadUop_io_uop_idx_valid = dec_io_isGemm ? tensorGemm_io_uop_idx_valid : tensorAlu_io_uop_idx_valid; // @[Compute.scala 120:22:@23286.4]
  assign loadUop_io_uop_idx_bits = dec_io_isGemm ? tensorGemm_io_uop_idx_bits : tensorAlu_io_uop_idx_bits; // @[Compute.scala 120:22:@23285.4]
  assign tensorAcc_clock = clock; // @[:@23204.4]
  assign tensorAcc_reset = reset; // @[:@23205.4]
  assign tensorAcc_io_start = _T_7083 & dec_io_isLoadAcc; // @[Compute.scala 123:22:@23290.4]
  assign tensorAcc_io_inst = inst_q_io_deq_bits; // @[Compute.scala 124:21:@23291.4]
  assign tensorAcc_io_baddr = io_acc_baddr; // @[Compute.scala 125:22:@23292.4]
  assign tensorAcc_io_vme_rd_cmd_ready = io_vme_rd_1_cmd_ready; // @[Compute.scala 128:16:@23321.4]
  assign tensorAcc_io_vme_rd_data_valid = io_vme_rd_1_data_valid; // @[Compute.scala 128:16:@23316.4]
  assign tensorAcc_io_vme_rd_data_bits = io_vme_rd_1_data_bits; // @[Compute.scala 128:16:@23315.4]
  assign tensorAcc_io_tensor_rd_idx_valid = dec_io_isGemm ? tensorGemm_io_acc_rd_idx_valid : tensorAlu_io_acc_rd_idx_valid; // @[Compute.scala 126:30:@23295.4]
  assign tensorAcc_io_tensor_rd_idx_bits = dec_io_isGemm ? tensorGemm_io_acc_rd_idx_bits : tensorAlu_io_acc_rd_idx_bits; // @[Compute.scala 126:30:@23294.4]
  assign tensorAcc_io_tensor_wr_valid = dec_io_isGemm ? tensorGemm_io_acc_wr_valid : tensorAlu_io_acc_wr_valid; // @[Compute.scala 127:26:@23314.4]
  assign tensorAcc_io_tensor_wr_bits_idx = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_idx : tensorAlu_io_acc_wr_bits_idx; // @[Compute.scala 127:26:@23313.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_0 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_0 : tensorAlu_io_acc_wr_bits_data_0_0; // @[Compute.scala 127:26:@23297.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_1 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_1 : tensorAlu_io_acc_wr_bits_data_0_1; // @[Compute.scala 127:26:@23298.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_2 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_2 : tensorAlu_io_acc_wr_bits_data_0_2; // @[Compute.scala 127:26:@23299.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_3 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_3 : tensorAlu_io_acc_wr_bits_data_0_3; // @[Compute.scala 127:26:@23300.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_4 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_4 : tensorAlu_io_acc_wr_bits_data_0_4; // @[Compute.scala 127:26:@23301.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_5 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_5 : tensorAlu_io_acc_wr_bits_data_0_5; // @[Compute.scala 127:26:@23302.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_6 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_6 : tensorAlu_io_acc_wr_bits_data_0_6; // @[Compute.scala 127:26:@23303.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_7 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_7 : tensorAlu_io_acc_wr_bits_data_0_7; // @[Compute.scala 127:26:@23304.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_8 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_8 : tensorAlu_io_acc_wr_bits_data_0_8; // @[Compute.scala 127:26:@23305.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_9 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_9 : tensorAlu_io_acc_wr_bits_data_0_9; // @[Compute.scala 127:26:@23306.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_10 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_10 : tensorAlu_io_acc_wr_bits_data_0_10; // @[Compute.scala 127:26:@23307.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_11 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_11 : tensorAlu_io_acc_wr_bits_data_0_11; // @[Compute.scala 127:26:@23308.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_12 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_12 : tensorAlu_io_acc_wr_bits_data_0_12; // @[Compute.scala 127:26:@23309.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_13 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_13 : tensorAlu_io_acc_wr_bits_data_0_13; // @[Compute.scala 127:26:@23310.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_14 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_14 : tensorAlu_io_acc_wr_bits_data_0_14; // @[Compute.scala 127:26:@23311.4]
  assign tensorAcc_io_tensor_wr_bits_data_0_15 = dec_io_isGemm ? tensorGemm_io_acc_wr_bits_data_0_15 : tensorAlu_io_acc_wr_bits_data_0_15; // @[Compute.scala 127:26:@23312.4]
  assign tensorGemm_clock = clock; // @[:@23207.4]
  assign tensorGemm_reset = reset; // @[:@23208.4]
  assign tensorGemm_io_start = _T_7083 & dec_io_isGemm; // @[Compute.scala 132:23:@23326.4]
  assign tensorGemm_io_inst = inst_q_io_deq_bits; // @[Compute.scala 133:22:@23327.4]
  assign tensorGemm_io_uop_data_valid = loadUop_io_uop_data_valid & dec_io_isGemm; // @[Compute.scala 134:32:@23329.4]
  assign tensorGemm_io_uop_data_bits_u2 = loadUop_io_uop_data_bits_u2; // @[Compute.scala 135:31:@23332.4]
  assign tensorGemm_io_uop_data_bits_u1 = loadUop_io_uop_data_bits_u1; // @[Compute.scala 135:31:@23331.4]
  assign tensorGemm_io_uop_data_bits_u0 = loadUop_io_uop_data_bits_u0; // @[Compute.scala 135:31:@23330.4]
  assign tensorGemm_io_inp_rd_data_valid = io_inp_rd_data_valid; // @[Compute.scala 136:21:@23367.4]
  assign tensorGemm_io_inp_rd_data_bits_0_0 = io_inp_rd_data_bits_0_0; // @[Compute.scala 136:21:@23351.4]
  assign tensorGemm_io_inp_rd_data_bits_0_1 = io_inp_rd_data_bits_0_1; // @[Compute.scala 136:21:@23352.4]
  assign tensorGemm_io_inp_rd_data_bits_0_2 = io_inp_rd_data_bits_0_2; // @[Compute.scala 136:21:@23353.4]
  assign tensorGemm_io_inp_rd_data_bits_0_3 = io_inp_rd_data_bits_0_3; // @[Compute.scala 136:21:@23354.4]
  assign tensorGemm_io_inp_rd_data_bits_0_4 = io_inp_rd_data_bits_0_4; // @[Compute.scala 136:21:@23355.4]
  assign tensorGemm_io_inp_rd_data_bits_0_5 = io_inp_rd_data_bits_0_5; // @[Compute.scala 136:21:@23356.4]
  assign tensorGemm_io_inp_rd_data_bits_0_6 = io_inp_rd_data_bits_0_6; // @[Compute.scala 136:21:@23357.4]
  assign tensorGemm_io_inp_rd_data_bits_0_7 = io_inp_rd_data_bits_0_7; // @[Compute.scala 136:21:@23358.4]
  assign tensorGemm_io_inp_rd_data_bits_0_8 = io_inp_rd_data_bits_0_8; // @[Compute.scala 136:21:@23359.4]
  assign tensorGemm_io_inp_rd_data_bits_0_9 = io_inp_rd_data_bits_0_9; // @[Compute.scala 136:21:@23360.4]
  assign tensorGemm_io_inp_rd_data_bits_0_10 = io_inp_rd_data_bits_0_10; // @[Compute.scala 136:21:@23361.4]
  assign tensorGemm_io_inp_rd_data_bits_0_11 = io_inp_rd_data_bits_0_11; // @[Compute.scala 136:21:@23362.4]
  assign tensorGemm_io_inp_rd_data_bits_0_12 = io_inp_rd_data_bits_0_12; // @[Compute.scala 136:21:@23363.4]
  assign tensorGemm_io_inp_rd_data_bits_0_13 = io_inp_rd_data_bits_0_13; // @[Compute.scala 136:21:@23364.4]
  assign tensorGemm_io_inp_rd_data_bits_0_14 = io_inp_rd_data_bits_0_14; // @[Compute.scala 136:21:@23365.4]
  assign tensorGemm_io_inp_rd_data_bits_0_15 = io_inp_rd_data_bits_0_15; // @[Compute.scala 136:21:@23366.4]
  assign tensorGemm_io_wgt_rd_data_valid = io_wgt_rd_data_valid; // @[Compute.scala 137:21:@23884.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_0 = io_wgt_rd_data_bits_0_0; // @[Compute.scala 137:21:@23628.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_1 = io_wgt_rd_data_bits_0_1; // @[Compute.scala 137:21:@23629.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_2 = io_wgt_rd_data_bits_0_2; // @[Compute.scala 137:21:@23630.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_3 = io_wgt_rd_data_bits_0_3; // @[Compute.scala 137:21:@23631.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_4 = io_wgt_rd_data_bits_0_4; // @[Compute.scala 137:21:@23632.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_5 = io_wgt_rd_data_bits_0_5; // @[Compute.scala 137:21:@23633.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_6 = io_wgt_rd_data_bits_0_6; // @[Compute.scala 137:21:@23634.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_7 = io_wgt_rd_data_bits_0_7; // @[Compute.scala 137:21:@23635.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_8 = io_wgt_rd_data_bits_0_8; // @[Compute.scala 137:21:@23636.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_9 = io_wgt_rd_data_bits_0_9; // @[Compute.scala 137:21:@23637.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_10 = io_wgt_rd_data_bits_0_10; // @[Compute.scala 137:21:@23638.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_11 = io_wgt_rd_data_bits_0_11; // @[Compute.scala 137:21:@23639.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_12 = io_wgt_rd_data_bits_0_12; // @[Compute.scala 137:21:@23640.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_13 = io_wgt_rd_data_bits_0_13; // @[Compute.scala 137:21:@23641.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_14 = io_wgt_rd_data_bits_0_14; // @[Compute.scala 137:21:@23642.4]
  assign tensorGemm_io_wgt_rd_data_bits_0_15 = io_wgt_rd_data_bits_0_15; // @[Compute.scala 137:21:@23643.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_0 = io_wgt_rd_data_bits_1_0; // @[Compute.scala 137:21:@23644.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_1 = io_wgt_rd_data_bits_1_1; // @[Compute.scala 137:21:@23645.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_2 = io_wgt_rd_data_bits_1_2; // @[Compute.scala 137:21:@23646.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_3 = io_wgt_rd_data_bits_1_3; // @[Compute.scala 137:21:@23647.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_4 = io_wgt_rd_data_bits_1_4; // @[Compute.scala 137:21:@23648.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_5 = io_wgt_rd_data_bits_1_5; // @[Compute.scala 137:21:@23649.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_6 = io_wgt_rd_data_bits_1_6; // @[Compute.scala 137:21:@23650.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_7 = io_wgt_rd_data_bits_1_7; // @[Compute.scala 137:21:@23651.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_8 = io_wgt_rd_data_bits_1_8; // @[Compute.scala 137:21:@23652.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_9 = io_wgt_rd_data_bits_1_9; // @[Compute.scala 137:21:@23653.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_10 = io_wgt_rd_data_bits_1_10; // @[Compute.scala 137:21:@23654.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_11 = io_wgt_rd_data_bits_1_11; // @[Compute.scala 137:21:@23655.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_12 = io_wgt_rd_data_bits_1_12; // @[Compute.scala 137:21:@23656.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_13 = io_wgt_rd_data_bits_1_13; // @[Compute.scala 137:21:@23657.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_14 = io_wgt_rd_data_bits_1_14; // @[Compute.scala 137:21:@23658.4]
  assign tensorGemm_io_wgt_rd_data_bits_1_15 = io_wgt_rd_data_bits_1_15; // @[Compute.scala 137:21:@23659.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_0 = io_wgt_rd_data_bits_2_0; // @[Compute.scala 137:21:@23660.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_1 = io_wgt_rd_data_bits_2_1; // @[Compute.scala 137:21:@23661.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_2 = io_wgt_rd_data_bits_2_2; // @[Compute.scala 137:21:@23662.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_3 = io_wgt_rd_data_bits_2_3; // @[Compute.scala 137:21:@23663.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_4 = io_wgt_rd_data_bits_2_4; // @[Compute.scala 137:21:@23664.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_5 = io_wgt_rd_data_bits_2_5; // @[Compute.scala 137:21:@23665.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_6 = io_wgt_rd_data_bits_2_6; // @[Compute.scala 137:21:@23666.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_7 = io_wgt_rd_data_bits_2_7; // @[Compute.scala 137:21:@23667.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_8 = io_wgt_rd_data_bits_2_8; // @[Compute.scala 137:21:@23668.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_9 = io_wgt_rd_data_bits_2_9; // @[Compute.scala 137:21:@23669.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_10 = io_wgt_rd_data_bits_2_10; // @[Compute.scala 137:21:@23670.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_11 = io_wgt_rd_data_bits_2_11; // @[Compute.scala 137:21:@23671.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_12 = io_wgt_rd_data_bits_2_12; // @[Compute.scala 137:21:@23672.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_13 = io_wgt_rd_data_bits_2_13; // @[Compute.scala 137:21:@23673.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_14 = io_wgt_rd_data_bits_2_14; // @[Compute.scala 137:21:@23674.4]
  assign tensorGemm_io_wgt_rd_data_bits_2_15 = io_wgt_rd_data_bits_2_15; // @[Compute.scala 137:21:@23675.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_0 = io_wgt_rd_data_bits_3_0; // @[Compute.scala 137:21:@23676.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_1 = io_wgt_rd_data_bits_3_1; // @[Compute.scala 137:21:@23677.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_2 = io_wgt_rd_data_bits_3_2; // @[Compute.scala 137:21:@23678.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_3 = io_wgt_rd_data_bits_3_3; // @[Compute.scala 137:21:@23679.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_4 = io_wgt_rd_data_bits_3_4; // @[Compute.scala 137:21:@23680.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_5 = io_wgt_rd_data_bits_3_5; // @[Compute.scala 137:21:@23681.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_6 = io_wgt_rd_data_bits_3_6; // @[Compute.scala 137:21:@23682.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_7 = io_wgt_rd_data_bits_3_7; // @[Compute.scala 137:21:@23683.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_8 = io_wgt_rd_data_bits_3_8; // @[Compute.scala 137:21:@23684.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_9 = io_wgt_rd_data_bits_3_9; // @[Compute.scala 137:21:@23685.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_10 = io_wgt_rd_data_bits_3_10; // @[Compute.scala 137:21:@23686.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_11 = io_wgt_rd_data_bits_3_11; // @[Compute.scala 137:21:@23687.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_12 = io_wgt_rd_data_bits_3_12; // @[Compute.scala 137:21:@23688.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_13 = io_wgt_rd_data_bits_3_13; // @[Compute.scala 137:21:@23689.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_14 = io_wgt_rd_data_bits_3_14; // @[Compute.scala 137:21:@23690.4]
  assign tensorGemm_io_wgt_rd_data_bits_3_15 = io_wgt_rd_data_bits_3_15; // @[Compute.scala 137:21:@23691.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_0 = io_wgt_rd_data_bits_4_0; // @[Compute.scala 137:21:@23692.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_1 = io_wgt_rd_data_bits_4_1; // @[Compute.scala 137:21:@23693.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_2 = io_wgt_rd_data_bits_4_2; // @[Compute.scala 137:21:@23694.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_3 = io_wgt_rd_data_bits_4_3; // @[Compute.scala 137:21:@23695.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_4 = io_wgt_rd_data_bits_4_4; // @[Compute.scala 137:21:@23696.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_5 = io_wgt_rd_data_bits_4_5; // @[Compute.scala 137:21:@23697.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_6 = io_wgt_rd_data_bits_4_6; // @[Compute.scala 137:21:@23698.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_7 = io_wgt_rd_data_bits_4_7; // @[Compute.scala 137:21:@23699.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_8 = io_wgt_rd_data_bits_4_8; // @[Compute.scala 137:21:@23700.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_9 = io_wgt_rd_data_bits_4_9; // @[Compute.scala 137:21:@23701.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_10 = io_wgt_rd_data_bits_4_10; // @[Compute.scala 137:21:@23702.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_11 = io_wgt_rd_data_bits_4_11; // @[Compute.scala 137:21:@23703.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_12 = io_wgt_rd_data_bits_4_12; // @[Compute.scala 137:21:@23704.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_13 = io_wgt_rd_data_bits_4_13; // @[Compute.scala 137:21:@23705.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_14 = io_wgt_rd_data_bits_4_14; // @[Compute.scala 137:21:@23706.4]
  assign tensorGemm_io_wgt_rd_data_bits_4_15 = io_wgt_rd_data_bits_4_15; // @[Compute.scala 137:21:@23707.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_0 = io_wgt_rd_data_bits_5_0; // @[Compute.scala 137:21:@23708.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_1 = io_wgt_rd_data_bits_5_1; // @[Compute.scala 137:21:@23709.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_2 = io_wgt_rd_data_bits_5_2; // @[Compute.scala 137:21:@23710.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_3 = io_wgt_rd_data_bits_5_3; // @[Compute.scala 137:21:@23711.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_4 = io_wgt_rd_data_bits_5_4; // @[Compute.scala 137:21:@23712.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_5 = io_wgt_rd_data_bits_5_5; // @[Compute.scala 137:21:@23713.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_6 = io_wgt_rd_data_bits_5_6; // @[Compute.scala 137:21:@23714.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_7 = io_wgt_rd_data_bits_5_7; // @[Compute.scala 137:21:@23715.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_8 = io_wgt_rd_data_bits_5_8; // @[Compute.scala 137:21:@23716.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_9 = io_wgt_rd_data_bits_5_9; // @[Compute.scala 137:21:@23717.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_10 = io_wgt_rd_data_bits_5_10; // @[Compute.scala 137:21:@23718.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_11 = io_wgt_rd_data_bits_5_11; // @[Compute.scala 137:21:@23719.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_12 = io_wgt_rd_data_bits_5_12; // @[Compute.scala 137:21:@23720.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_13 = io_wgt_rd_data_bits_5_13; // @[Compute.scala 137:21:@23721.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_14 = io_wgt_rd_data_bits_5_14; // @[Compute.scala 137:21:@23722.4]
  assign tensorGemm_io_wgt_rd_data_bits_5_15 = io_wgt_rd_data_bits_5_15; // @[Compute.scala 137:21:@23723.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_0 = io_wgt_rd_data_bits_6_0; // @[Compute.scala 137:21:@23724.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_1 = io_wgt_rd_data_bits_6_1; // @[Compute.scala 137:21:@23725.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_2 = io_wgt_rd_data_bits_6_2; // @[Compute.scala 137:21:@23726.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_3 = io_wgt_rd_data_bits_6_3; // @[Compute.scala 137:21:@23727.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_4 = io_wgt_rd_data_bits_6_4; // @[Compute.scala 137:21:@23728.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_5 = io_wgt_rd_data_bits_6_5; // @[Compute.scala 137:21:@23729.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_6 = io_wgt_rd_data_bits_6_6; // @[Compute.scala 137:21:@23730.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_7 = io_wgt_rd_data_bits_6_7; // @[Compute.scala 137:21:@23731.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_8 = io_wgt_rd_data_bits_6_8; // @[Compute.scala 137:21:@23732.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_9 = io_wgt_rd_data_bits_6_9; // @[Compute.scala 137:21:@23733.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_10 = io_wgt_rd_data_bits_6_10; // @[Compute.scala 137:21:@23734.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_11 = io_wgt_rd_data_bits_6_11; // @[Compute.scala 137:21:@23735.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_12 = io_wgt_rd_data_bits_6_12; // @[Compute.scala 137:21:@23736.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_13 = io_wgt_rd_data_bits_6_13; // @[Compute.scala 137:21:@23737.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_14 = io_wgt_rd_data_bits_6_14; // @[Compute.scala 137:21:@23738.4]
  assign tensorGemm_io_wgt_rd_data_bits_6_15 = io_wgt_rd_data_bits_6_15; // @[Compute.scala 137:21:@23739.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_0 = io_wgt_rd_data_bits_7_0; // @[Compute.scala 137:21:@23740.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_1 = io_wgt_rd_data_bits_7_1; // @[Compute.scala 137:21:@23741.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_2 = io_wgt_rd_data_bits_7_2; // @[Compute.scala 137:21:@23742.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_3 = io_wgt_rd_data_bits_7_3; // @[Compute.scala 137:21:@23743.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_4 = io_wgt_rd_data_bits_7_4; // @[Compute.scala 137:21:@23744.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_5 = io_wgt_rd_data_bits_7_5; // @[Compute.scala 137:21:@23745.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_6 = io_wgt_rd_data_bits_7_6; // @[Compute.scala 137:21:@23746.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_7 = io_wgt_rd_data_bits_7_7; // @[Compute.scala 137:21:@23747.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_8 = io_wgt_rd_data_bits_7_8; // @[Compute.scala 137:21:@23748.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_9 = io_wgt_rd_data_bits_7_9; // @[Compute.scala 137:21:@23749.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_10 = io_wgt_rd_data_bits_7_10; // @[Compute.scala 137:21:@23750.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_11 = io_wgt_rd_data_bits_7_11; // @[Compute.scala 137:21:@23751.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_12 = io_wgt_rd_data_bits_7_12; // @[Compute.scala 137:21:@23752.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_13 = io_wgt_rd_data_bits_7_13; // @[Compute.scala 137:21:@23753.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_14 = io_wgt_rd_data_bits_7_14; // @[Compute.scala 137:21:@23754.4]
  assign tensorGemm_io_wgt_rd_data_bits_7_15 = io_wgt_rd_data_bits_7_15; // @[Compute.scala 137:21:@23755.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_0 = io_wgt_rd_data_bits_8_0; // @[Compute.scala 137:21:@23756.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_1 = io_wgt_rd_data_bits_8_1; // @[Compute.scala 137:21:@23757.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_2 = io_wgt_rd_data_bits_8_2; // @[Compute.scala 137:21:@23758.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_3 = io_wgt_rd_data_bits_8_3; // @[Compute.scala 137:21:@23759.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_4 = io_wgt_rd_data_bits_8_4; // @[Compute.scala 137:21:@23760.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_5 = io_wgt_rd_data_bits_8_5; // @[Compute.scala 137:21:@23761.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_6 = io_wgt_rd_data_bits_8_6; // @[Compute.scala 137:21:@23762.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_7 = io_wgt_rd_data_bits_8_7; // @[Compute.scala 137:21:@23763.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_8 = io_wgt_rd_data_bits_8_8; // @[Compute.scala 137:21:@23764.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_9 = io_wgt_rd_data_bits_8_9; // @[Compute.scala 137:21:@23765.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_10 = io_wgt_rd_data_bits_8_10; // @[Compute.scala 137:21:@23766.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_11 = io_wgt_rd_data_bits_8_11; // @[Compute.scala 137:21:@23767.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_12 = io_wgt_rd_data_bits_8_12; // @[Compute.scala 137:21:@23768.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_13 = io_wgt_rd_data_bits_8_13; // @[Compute.scala 137:21:@23769.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_14 = io_wgt_rd_data_bits_8_14; // @[Compute.scala 137:21:@23770.4]
  assign tensorGemm_io_wgt_rd_data_bits_8_15 = io_wgt_rd_data_bits_8_15; // @[Compute.scala 137:21:@23771.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_0 = io_wgt_rd_data_bits_9_0; // @[Compute.scala 137:21:@23772.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_1 = io_wgt_rd_data_bits_9_1; // @[Compute.scala 137:21:@23773.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_2 = io_wgt_rd_data_bits_9_2; // @[Compute.scala 137:21:@23774.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_3 = io_wgt_rd_data_bits_9_3; // @[Compute.scala 137:21:@23775.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_4 = io_wgt_rd_data_bits_9_4; // @[Compute.scala 137:21:@23776.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_5 = io_wgt_rd_data_bits_9_5; // @[Compute.scala 137:21:@23777.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_6 = io_wgt_rd_data_bits_9_6; // @[Compute.scala 137:21:@23778.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_7 = io_wgt_rd_data_bits_9_7; // @[Compute.scala 137:21:@23779.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_8 = io_wgt_rd_data_bits_9_8; // @[Compute.scala 137:21:@23780.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_9 = io_wgt_rd_data_bits_9_9; // @[Compute.scala 137:21:@23781.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_10 = io_wgt_rd_data_bits_9_10; // @[Compute.scala 137:21:@23782.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_11 = io_wgt_rd_data_bits_9_11; // @[Compute.scala 137:21:@23783.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_12 = io_wgt_rd_data_bits_9_12; // @[Compute.scala 137:21:@23784.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_13 = io_wgt_rd_data_bits_9_13; // @[Compute.scala 137:21:@23785.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_14 = io_wgt_rd_data_bits_9_14; // @[Compute.scala 137:21:@23786.4]
  assign tensorGemm_io_wgt_rd_data_bits_9_15 = io_wgt_rd_data_bits_9_15; // @[Compute.scala 137:21:@23787.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_0 = io_wgt_rd_data_bits_10_0; // @[Compute.scala 137:21:@23788.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_1 = io_wgt_rd_data_bits_10_1; // @[Compute.scala 137:21:@23789.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_2 = io_wgt_rd_data_bits_10_2; // @[Compute.scala 137:21:@23790.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_3 = io_wgt_rd_data_bits_10_3; // @[Compute.scala 137:21:@23791.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_4 = io_wgt_rd_data_bits_10_4; // @[Compute.scala 137:21:@23792.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_5 = io_wgt_rd_data_bits_10_5; // @[Compute.scala 137:21:@23793.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_6 = io_wgt_rd_data_bits_10_6; // @[Compute.scala 137:21:@23794.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_7 = io_wgt_rd_data_bits_10_7; // @[Compute.scala 137:21:@23795.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_8 = io_wgt_rd_data_bits_10_8; // @[Compute.scala 137:21:@23796.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_9 = io_wgt_rd_data_bits_10_9; // @[Compute.scala 137:21:@23797.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_10 = io_wgt_rd_data_bits_10_10; // @[Compute.scala 137:21:@23798.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_11 = io_wgt_rd_data_bits_10_11; // @[Compute.scala 137:21:@23799.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_12 = io_wgt_rd_data_bits_10_12; // @[Compute.scala 137:21:@23800.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_13 = io_wgt_rd_data_bits_10_13; // @[Compute.scala 137:21:@23801.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_14 = io_wgt_rd_data_bits_10_14; // @[Compute.scala 137:21:@23802.4]
  assign tensorGemm_io_wgt_rd_data_bits_10_15 = io_wgt_rd_data_bits_10_15; // @[Compute.scala 137:21:@23803.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_0 = io_wgt_rd_data_bits_11_0; // @[Compute.scala 137:21:@23804.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_1 = io_wgt_rd_data_bits_11_1; // @[Compute.scala 137:21:@23805.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_2 = io_wgt_rd_data_bits_11_2; // @[Compute.scala 137:21:@23806.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_3 = io_wgt_rd_data_bits_11_3; // @[Compute.scala 137:21:@23807.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_4 = io_wgt_rd_data_bits_11_4; // @[Compute.scala 137:21:@23808.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_5 = io_wgt_rd_data_bits_11_5; // @[Compute.scala 137:21:@23809.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_6 = io_wgt_rd_data_bits_11_6; // @[Compute.scala 137:21:@23810.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_7 = io_wgt_rd_data_bits_11_7; // @[Compute.scala 137:21:@23811.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_8 = io_wgt_rd_data_bits_11_8; // @[Compute.scala 137:21:@23812.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_9 = io_wgt_rd_data_bits_11_9; // @[Compute.scala 137:21:@23813.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_10 = io_wgt_rd_data_bits_11_10; // @[Compute.scala 137:21:@23814.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_11 = io_wgt_rd_data_bits_11_11; // @[Compute.scala 137:21:@23815.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_12 = io_wgt_rd_data_bits_11_12; // @[Compute.scala 137:21:@23816.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_13 = io_wgt_rd_data_bits_11_13; // @[Compute.scala 137:21:@23817.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_14 = io_wgt_rd_data_bits_11_14; // @[Compute.scala 137:21:@23818.4]
  assign tensorGemm_io_wgt_rd_data_bits_11_15 = io_wgt_rd_data_bits_11_15; // @[Compute.scala 137:21:@23819.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_0 = io_wgt_rd_data_bits_12_0; // @[Compute.scala 137:21:@23820.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_1 = io_wgt_rd_data_bits_12_1; // @[Compute.scala 137:21:@23821.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_2 = io_wgt_rd_data_bits_12_2; // @[Compute.scala 137:21:@23822.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_3 = io_wgt_rd_data_bits_12_3; // @[Compute.scala 137:21:@23823.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_4 = io_wgt_rd_data_bits_12_4; // @[Compute.scala 137:21:@23824.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_5 = io_wgt_rd_data_bits_12_5; // @[Compute.scala 137:21:@23825.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_6 = io_wgt_rd_data_bits_12_6; // @[Compute.scala 137:21:@23826.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_7 = io_wgt_rd_data_bits_12_7; // @[Compute.scala 137:21:@23827.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_8 = io_wgt_rd_data_bits_12_8; // @[Compute.scala 137:21:@23828.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_9 = io_wgt_rd_data_bits_12_9; // @[Compute.scala 137:21:@23829.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_10 = io_wgt_rd_data_bits_12_10; // @[Compute.scala 137:21:@23830.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_11 = io_wgt_rd_data_bits_12_11; // @[Compute.scala 137:21:@23831.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_12 = io_wgt_rd_data_bits_12_12; // @[Compute.scala 137:21:@23832.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_13 = io_wgt_rd_data_bits_12_13; // @[Compute.scala 137:21:@23833.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_14 = io_wgt_rd_data_bits_12_14; // @[Compute.scala 137:21:@23834.4]
  assign tensorGemm_io_wgt_rd_data_bits_12_15 = io_wgt_rd_data_bits_12_15; // @[Compute.scala 137:21:@23835.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_0 = io_wgt_rd_data_bits_13_0; // @[Compute.scala 137:21:@23836.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_1 = io_wgt_rd_data_bits_13_1; // @[Compute.scala 137:21:@23837.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_2 = io_wgt_rd_data_bits_13_2; // @[Compute.scala 137:21:@23838.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_3 = io_wgt_rd_data_bits_13_3; // @[Compute.scala 137:21:@23839.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_4 = io_wgt_rd_data_bits_13_4; // @[Compute.scala 137:21:@23840.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_5 = io_wgt_rd_data_bits_13_5; // @[Compute.scala 137:21:@23841.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_6 = io_wgt_rd_data_bits_13_6; // @[Compute.scala 137:21:@23842.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_7 = io_wgt_rd_data_bits_13_7; // @[Compute.scala 137:21:@23843.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_8 = io_wgt_rd_data_bits_13_8; // @[Compute.scala 137:21:@23844.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_9 = io_wgt_rd_data_bits_13_9; // @[Compute.scala 137:21:@23845.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_10 = io_wgt_rd_data_bits_13_10; // @[Compute.scala 137:21:@23846.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_11 = io_wgt_rd_data_bits_13_11; // @[Compute.scala 137:21:@23847.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_12 = io_wgt_rd_data_bits_13_12; // @[Compute.scala 137:21:@23848.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_13 = io_wgt_rd_data_bits_13_13; // @[Compute.scala 137:21:@23849.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_14 = io_wgt_rd_data_bits_13_14; // @[Compute.scala 137:21:@23850.4]
  assign tensorGemm_io_wgt_rd_data_bits_13_15 = io_wgt_rd_data_bits_13_15; // @[Compute.scala 137:21:@23851.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_0 = io_wgt_rd_data_bits_14_0; // @[Compute.scala 137:21:@23852.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_1 = io_wgt_rd_data_bits_14_1; // @[Compute.scala 137:21:@23853.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_2 = io_wgt_rd_data_bits_14_2; // @[Compute.scala 137:21:@23854.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_3 = io_wgt_rd_data_bits_14_3; // @[Compute.scala 137:21:@23855.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_4 = io_wgt_rd_data_bits_14_4; // @[Compute.scala 137:21:@23856.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_5 = io_wgt_rd_data_bits_14_5; // @[Compute.scala 137:21:@23857.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_6 = io_wgt_rd_data_bits_14_6; // @[Compute.scala 137:21:@23858.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_7 = io_wgt_rd_data_bits_14_7; // @[Compute.scala 137:21:@23859.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_8 = io_wgt_rd_data_bits_14_8; // @[Compute.scala 137:21:@23860.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_9 = io_wgt_rd_data_bits_14_9; // @[Compute.scala 137:21:@23861.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_10 = io_wgt_rd_data_bits_14_10; // @[Compute.scala 137:21:@23862.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_11 = io_wgt_rd_data_bits_14_11; // @[Compute.scala 137:21:@23863.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_12 = io_wgt_rd_data_bits_14_12; // @[Compute.scala 137:21:@23864.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_13 = io_wgt_rd_data_bits_14_13; // @[Compute.scala 137:21:@23865.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_14 = io_wgt_rd_data_bits_14_14; // @[Compute.scala 137:21:@23866.4]
  assign tensorGemm_io_wgt_rd_data_bits_14_15 = io_wgt_rd_data_bits_14_15; // @[Compute.scala 137:21:@23867.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_0 = io_wgt_rd_data_bits_15_0; // @[Compute.scala 137:21:@23868.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_1 = io_wgt_rd_data_bits_15_1; // @[Compute.scala 137:21:@23869.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_2 = io_wgt_rd_data_bits_15_2; // @[Compute.scala 137:21:@23870.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_3 = io_wgt_rd_data_bits_15_3; // @[Compute.scala 137:21:@23871.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_4 = io_wgt_rd_data_bits_15_4; // @[Compute.scala 137:21:@23872.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_5 = io_wgt_rd_data_bits_15_5; // @[Compute.scala 137:21:@23873.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_6 = io_wgt_rd_data_bits_15_6; // @[Compute.scala 137:21:@23874.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_7 = io_wgt_rd_data_bits_15_7; // @[Compute.scala 137:21:@23875.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_8 = io_wgt_rd_data_bits_15_8; // @[Compute.scala 137:21:@23876.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_9 = io_wgt_rd_data_bits_15_9; // @[Compute.scala 137:21:@23877.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_10 = io_wgt_rd_data_bits_15_10; // @[Compute.scala 137:21:@23878.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_11 = io_wgt_rd_data_bits_15_11; // @[Compute.scala 137:21:@23879.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_12 = io_wgt_rd_data_bits_15_12; // @[Compute.scala 137:21:@23880.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_13 = io_wgt_rd_data_bits_15_13; // @[Compute.scala 137:21:@23881.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_14 = io_wgt_rd_data_bits_15_14; // @[Compute.scala 137:21:@23882.4]
  assign tensorGemm_io_wgt_rd_data_bits_15_15 = io_wgt_rd_data_bits_15_15; // @[Compute.scala 137:21:@23883.4]
  assign tensorGemm_io_acc_rd_data_valid = tensorAcc_io_tensor_rd_data_valid & dec_io_isGemm; // @[Compute.scala 138:35:@23888.4]
  assign tensorGemm_io_acc_rd_data_bits_0_0 = tensorAcc_io_tensor_rd_data_bits_0_0; // @[Compute.scala 139:34:@23889.4]
  assign tensorGemm_io_acc_rd_data_bits_0_1 = tensorAcc_io_tensor_rd_data_bits_0_1; // @[Compute.scala 139:34:@23890.4]
  assign tensorGemm_io_acc_rd_data_bits_0_2 = tensorAcc_io_tensor_rd_data_bits_0_2; // @[Compute.scala 139:34:@23891.4]
  assign tensorGemm_io_acc_rd_data_bits_0_3 = tensorAcc_io_tensor_rd_data_bits_0_3; // @[Compute.scala 139:34:@23892.4]
  assign tensorGemm_io_acc_rd_data_bits_0_4 = tensorAcc_io_tensor_rd_data_bits_0_4; // @[Compute.scala 139:34:@23893.4]
  assign tensorGemm_io_acc_rd_data_bits_0_5 = tensorAcc_io_tensor_rd_data_bits_0_5; // @[Compute.scala 139:34:@23894.4]
  assign tensorGemm_io_acc_rd_data_bits_0_6 = tensorAcc_io_tensor_rd_data_bits_0_6; // @[Compute.scala 139:34:@23895.4]
  assign tensorGemm_io_acc_rd_data_bits_0_7 = tensorAcc_io_tensor_rd_data_bits_0_7; // @[Compute.scala 139:34:@23896.4]
  assign tensorGemm_io_acc_rd_data_bits_0_8 = tensorAcc_io_tensor_rd_data_bits_0_8; // @[Compute.scala 139:34:@23897.4]
  assign tensorGemm_io_acc_rd_data_bits_0_9 = tensorAcc_io_tensor_rd_data_bits_0_9; // @[Compute.scala 139:34:@23898.4]
  assign tensorGemm_io_acc_rd_data_bits_0_10 = tensorAcc_io_tensor_rd_data_bits_0_10; // @[Compute.scala 139:34:@23899.4]
  assign tensorGemm_io_acc_rd_data_bits_0_11 = tensorAcc_io_tensor_rd_data_bits_0_11; // @[Compute.scala 139:34:@23900.4]
  assign tensorGemm_io_acc_rd_data_bits_0_12 = tensorAcc_io_tensor_rd_data_bits_0_12; // @[Compute.scala 139:34:@23901.4]
  assign tensorGemm_io_acc_rd_data_bits_0_13 = tensorAcc_io_tensor_rd_data_bits_0_13; // @[Compute.scala 139:34:@23902.4]
  assign tensorGemm_io_acc_rd_data_bits_0_14 = tensorAcc_io_tensor_rd_data_bits_0_14; // @[Compute.scala 139:34:@23903.4]
  assign tensorGemm_io_acc_rd_data_bits_0_15 = tensorAcc_io_tensor_rd_data_bits_0_15; // @[Compute.scala 139:34:@23904.4]
  assign tensorAlu_clock = clock; // @[:@23210.4]
  assign tensorAlu_reset = reset; // @[:@23211.4]
  assign tensorAlu_io_start = _T_7083 & dec_io_isAlu; // @[Compute.scala 144:22:@23926.4]
  assign tensorAlu_io_inst = inst_q_io_deq_bits; // @[Compute.scala 145:21:@23927.4]
  assign tensorAlu_io_uop_data_valid = loadUop_io_uop_data_valid & dec_io_isAlu; // @[Compute.scala 146:31:@23929.4]
  assign tensorAlu_io_uop_data_bits_u1 = loadUop_io_uop_data_bits_u1; // @[Compute.scala 147:30:@23931.4]
  assign tensorAlu_io_uop_data_bits_u0 = loadUop_io_uop_data_bits_u0; // @[Compute.scala 147:30:@23930.4]
  assign tensorAlu_io_acc_rd_data_valid = tensorAcc_io_tensor_rd_data_valid & dec_io_isAlu; // @[Compute.scala 148:34:@23934.4]
  assign tensorAlu_io_acc_rd_data_bits_0_0 = tensorAcc_io_tensor_rd_data_bits_0_0; // @[Compute.scala 149:33:@23935.4]
  assign tensorAlu_io_acc_rd_data_bits_0_1 = tensorAcc_io_tensor_rd_data_bits_0_1; // @[Compute.scala 149:33:@23936.4]
  assign tensorAlu_io_acc_rd_data_bits_0_2 = tensorAcc_io_tensor_rd_data_bits_0_2; // @[Compute.scala 149:33:@23937.4]
  assign tensorAlu_io_acc_rd_data_bits_0_3 = tensorAcc_io_tensor_rd_data_bits_0_3; // @[Compute.scala 149:33:@23938.4]
  assign tensorAlu_io_acc_rd_data_bits_0_4 = tensorAcc_io_tensor_rd_data_bits_0_4; // @[Compute.scala 149:33:@23939.4]
  assign tensorAlu_io_acc_rd_data_bits_0_5 = tensorAcc_io_tensor_rd_data_bits_0_5; // @[Compute.scala 149:33:@23940.4]
  assign tensorAlu_io_acc_rd_data_bits_0_6 = tensorAcc_io_tensor_rd_data_bits_0_6; // @[Compute.scala 149:33:@23941.4]
  assign tensorAlu_io_acc_rd_data_bits_0_7 = tensorAcc_io_tensor_rd_data_bits_0_7; // @[Compute.scala 149:33:@23942.4]
  assign tensorAlu_io_acc_rd_data_bits_0_8 = tensorAcc_io_tensor_rd_data_bits_0_8; // @[Compute.scala 149:33:@23943.4]
  assign tensorAlu_io_acc_rd_data_bits_0_9 = tensorAcc_io_tensor_rd_data_bits_0_9; // @[Compute.scala 149:33:@23944.4]
  assign tensorAlu_io_acc_rd_data_bits_0_10 = tensorAcc_io_tensor_rd_data_bits_0_10; // @[Compute.scala 149:33:@23945.4]
  assign tensorAlu_io_acc_rd_data_bits_0_11 = tensorAcc_io_tensor_rd_data_bits_0_11; // @[Compute.scala 149:33:@23946.4]
  assign tensorAlu_io_acc_rd_data_bits_0_12 = tensorAcc_io_tensor_rd_data_bits_0_12; // @[Compute.scala 149:33:@23947.4]
  assign tensorAlu_io_acc_rd_data_bits_0_13 = tensorAcc_io_tensor_rd_data_bits_0_13; // @[Compute.scala 149:33:@23948.4]
  assign tensorAlu_io_acc_rd_data_bits_0_14 = tensorAcc_io_tensor_rd_data_bits_0_14; // @[Compute.scala 149:33:@23949.4]
  assign tensorAlu_io_acc_rd_data_bits_0_15 = tensorAcc_io_tensor_rd_data_bits_0_15; // @[Compute.scala 149:33:@23950.4]
  assign inst_q_clock = clock; // @[:@23213.4]
  assign inst_q_reset = reset; // @[:@23214.4]
  assign inst_q_io_enq_valid = io_inst_valid; // @[Compute.scala 112:17:@23264.4]
  assign inst_q_io_enq_bits = io_inst_bits; // @[Compute.scala 112:17:@23263.4]
  assign inst_q_io_deq_ready = _T_7079 | _T_7080; // @[Compute.scala 113:23:@23270.4]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Compute.scala 65:15:@23218.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_7073) begin
        if (start) begin
          if (dec_io_isSync) begin
            state <= 2'h1;
          end else begin
            if (_T_7075) begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_7076) begin
          state <= 2'h0;
        end else begin
          if (_T_7077) begin
            if (done) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module StoreDecode( // @[:@24097.2]
  input  [127:0] io_inst, // @[:@24100.4]
  output         io_push_prev, // @[:@24100.4]
  output         io_pop_prev, // @[:@24100.4]
  output         io_isStore, // @[:@24100.4]
  output         io_isSync // @[:@24100.4]
);
  wire [15:0] dec_xsize; // @[Decode.scala 225:29:@24125.4]
  wire [127:0] _T_37; // @[Decode.scala 228:25:@24139.4]
  wire  _T_38; // @[Decode.scala 228:25:@24140.4]
  wire  _T_40; // @[Decode.scala 228:46:@24141.4]
  wire  _T_47; // @[Decode.scala 229:45:@24146.4]
  assign dec_xsize = io_inst[95:80]; // @[Decode.scala 225:29:@24125.4]
  assign _T_37 = io_inst & 128'h7; // @[Decode.scala 228:25:@24139.4]
  assign _T_38 = 128'h1 == _T_37; // @[Decode.scala 228:25:@24140.4]
  assign _T_40 = dec_xsize != 16'h0; // @[Decode.scala 228:46:@24141.4]
  assign _T_47 = dec_xsize == 16'h0; // @[Decode.scala 229:45:@24146.4]
  assign io_push_prev = io_inst[5]; // @[Decode.scala 226:16:@24137.4]
  assign io_pop_prev = io_inst[3]; // @[Decode.scala 227:15:@24138.4]
  assign io_isStore = _T_38 & _T_40; // @[Decode.scala 228:14:@24143.4]
  assign io_isSync = _T_38 & _T_47; // @[Decode.scala 229:13:@24148.4]
endmodule
module TensorStore( // @[:@24150.2]
  input          clock, // @[:@24151.4]
  input          reset, // @[:@24152.4]
  input          io_start, // @[:@24153.4]
  output         io_done, // @[:@24153.4]
  input  [127:0] io_inst, // @[:@24153.4]
  input  [31:0]  io_baddr, // @[:@24153.4]
  input          io_vme_wr_cmd_ready, // @[:@24153.4]
  output         io_vme_wr_cmd_valid, // @[:@24153.4]
  output [31:0]  io_vme_wr_cmd_bits_addr, // @[:@24153.4]
  output [7:0]   io_vme_wr_cmd_bits_len, // @[:@24153.4]
  input          io_vme_wr_data_ready, // @[:@24153.4]
  output         io_vme_wr_data_valid, // @[:@24153.4]
  output [63:0]  io_vme_wr_data_bits, // @[:@24153.4]
  input          io_vme_wr_ack, // @[:@24153.4]
  input          io_tensor_wr_valid, // @[:@24153.4]
  input  [10:0]  io_tensor_wr_bits_idx, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_0, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_1, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_2, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_3, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_4, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_5, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_6, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_7, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_8, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_9, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_10, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_11, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_12, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_13, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_14, // @[:@24153.4]
  input  [7:0]   io_tensor_wr_bits_data_0_15 // @[:@24153.4]
);
  reg [63:0] tensorFile_0_0 [0:2047]; // @[TensorStore.scala 152:16:@24395.4]
  reg [63:0] _RAND_0;
  wire [63:0] tensorFile_0_0__T_914_data; // @[TensorStore.scala 152:16:@24395.4]
  wire [10:0] tensorFile_0_0__T_914_addr; // @[TensorStore.scala 152:16:@24395.4]
  wire [63:0] tensorFile_0_0__T_836_data; // @[TensorStore.scala 152:16:@24395.4]
  wire [10:0] tensorFile_0_0__T_836_addr; // @[TensorStore.scala 152:16:@24395.4]
  wire  tensorFile_0_0__T_836_mask; // @[TensorStore.scala 152:16:@24395.4]
  wire  tensorFile_0_0__T_836_en; // @[TensorStore.scala 152:16:@24395.4]
  reg [63:0] tensorFile_0_1 [0:2047]; // @[TensorStore.scala 152:16:@24395.4]
  reg [63:0] _RAND_1;
  wire [63:0] tensorFile_0_1__T_914_data; // @[TensorStore.scala 152:16:@24395.4]
  wire [10:0] tensorFile_0_1__T_914_addr; // @[TensorStore.scala 152:16:@24395.4]
  wire [63:0] tensorFile_0_1__T_836_data; // @[TensorStore.scala 152:16:@24395.4]
  wire [10:0] tensorFile_0_1__T_836_addr; // @[TensorStore.scala 152:16:@24395.4]
  wire  tensorFile_0_1__T_836_mask; // @[TensorStore.scala 152:16:@24395.4]
  wire  tensorFile_0_1__T_836_en; // @[TensorStore.scala 152:16:@24395.4]
  wire [15:0] dec_sram_offset; // @[TensorStore.scala 51:29:@24170.4]
  wire [31:0] dec_dram_offset; // @[TensorStore.scala 51:29:@24172.4]
  wire [15:0] dec_ysize; // @[TensorStore.scala 51:29:@24176.4]
  wire [15:0] dec_xsize; // @[TensorStore.scala 51:29:@24178.4]
  wire [15:0] dec_xstride; // @[TensorStore.scala 51:29:@24180.4]
  reg [31:0] waddr_cur; // @[TensorStore.scala 52:22:@24190.4]
  reg [31:0] _RAND_2;
  reg [31:0] waddr_nxt; // @[TensorStore.scala 53:22:@24191.4]
  reg [31:0] _RAND_3;
  reg [7:0] xcnt; // @[TensorStore.scala 54:17:@24192.4]
  reg [31:0] _RAND_4;
  reg [7:0] xlen; // @[TensorStore.scala 55:17:@24193.4]
  reg [31:0] _RAND_5;
  reg [15:0] xrem; // @[TensorStore.scala 56:17:@24194.4]
  reg [31:0] _RAND_6;
  wire [16:0] _GEN_96; // @[TensorStore.scala 57:26:@24195.4]
  wire [16:0] _T_610; // @[TensorStore.scala 57:26:@24195.4]
  wire [17:0] _T_612; // @[TensorStore.scala 57:67:@24196.4]
  wire [17:0] _T_613; // @[TensorStore.scala 57:67:@24197.4]
  wire [16:0] xsize; // @[TensorStore.scala 57:67:@24198.4]
  reg [15:0] ycnt; // @[TensorStore.scala 60:17:@24199.4]
  reg [31:0] _RAND_7;
  reg [7:0] tag; // @[TensorStore.scala 62:16:@24200.4]
  reg [31:0] _RAND_8;
  reg [7:0] set; // @[TensorStore.scala 63:16:@24201.4]
  reg [31:0] _RAND_9;
  reg [31:0] xfer_bytes; // @[TensorStore.scala 65:23:@24202.4]
  reg [31:0] _RAND_10;
  wire [19:0] _GEN_97; // @[TensorStore.scala 66:35:@24203.4]
  wire [19:0] xstride_bytes; // @[TensorStore.scala 66:35:@24203.4]
  wire [35:0] _GEN_98; // @[TensorStore.scala 71:66:@24268.4]
  wire [35:0] _T_718; // @[TensorStore.scala 71:66:@24268.4]
  wire [35:0] _T_719; // @[TensorStore.scala 71:47:@24269.4]
  wire [35:0] _GEN_99; // @[TensorStore.scala 71:33:@24270.4]
  wire [35:0] xfer_init_addr; // @[TensorStore.scala 71:33:@24270.4]
  wire [32:0] _T_720; // @[TensorStore.scala 72:35:@24271.4]
  wire [31:0] xfer_split_addr; // @[TensorStore.scala 72:35:@24272.4]
  wire [31:0] _GEN_100; // @[TensorStore.scala 73:36:@24273.4]
  wire [32:0] _T_721; // @[TensorStore.scala 73:36:@24273.4]
  wire [31:0] xfer_stride_addr; // @[TensorStore.scala 73:36:@24274.4]
  wire [35:0] _GEN_15; // @[TensorStore.scala 75:55:@24275.4]
  wire [11:0] _T_722; // @[TensorStore.scala 75:55:@24275.4]
  wire [12:0] _T_723; // @[TensorStore.scala 75:38:@24276.4]
  wire [12:0] _T_724; // @[TensorStore.scala 75:38:@24277.4]
  wire [11:0] xfer_init_bytes; // @[TensorStore.scala 75:38:@24278.4]
  wire [8:0] xfer_init_pulses; // @[TensorStore.scala 76:43:@24279.4]
  wire [31:0] _GEN_16; // @[TensorStore.scala 77:56:@24280.4]
  wire [11:0] _T_725; // @[TensorStore.scala 77:56:@24280.4]
  wire [12:0] _T_726; // @[TensorStore.scala 77:38:@24281.4]
  wire [12:0] _T_727; // @[TensorStore.scala 77:38:@24282.4]
  wire [11:0] xfer_split_bytes; // @[TensorStore.scala 77:38:@24283.4]
  wire [8:0] xfer_split_pulses; // @[TensorStore.scala 78:44:@24284.4]
  wire [31:0] _GEN_43; // @[TensorStore.scala 79:57:@24285.4]
  wire [11:0] _T_728; // @[TensorStore.scala 79:57:@24285.4]
  wire [12:0] _T_729; // @[TensorStore.scala 79:38:@24286.4]
  wire [12:0] _T_730; // @[TensorStore.scala 79:38:@24287.4]
  wire [11:0] xfer_stride_bytes; // @[TensorStore.scala 79:38:@24288.4]
  wire [8:0] xfer_stride_pulses; // @[TensorStore.scala 80:45:@24289.4]
  reg [2:0] state; // @[TensorStore.scala 83:22:@24290.4]
  reg [31:0] _RAND_11;
  wire  _T_732; // @[Conditional.scala 37:30:@24291.4]
  wire [16:0] _GEN_101; // @[TensorStore.scala 91:21:@24296.8]
  wire  _T_733; // @[TensorStore.scala 91:21:@24296.8]
  wire [9:0] _T_736; // @[TensorStore.scala 95:36:@24302.10]
  wire [9:0] _T_737; // @[TensorStore.scala 95:36:@24303.10]
  wire [8:0] _T_738; // @[TensorStore.scala 95:36:@24304.10]
  wire [17:0] _T_739; // @[TensorStore.scala 96:25:@24306.10]
  wire [17:0] _T_740; // @[TensorStore.scala 96:25:@24307.10]
  wire [16:0] _T_741; // @[TensorStore.scala 96:25:@24308.10]
  wire [16:0] _GEN_0; // @[TensorStore.scala 91:41:@24297.8]
  wire [16:0] _GEN_1; // @[TensorStore.scala 91:41:@24297.8]
  wire [2:0] _GEN_2; // @[TensorStore.scala 89:23:@24294.6]
  wire [16:0] _GEN_3; // @[TensorStore.scala 89:23:@24294.6]
  wire [16:0] _GEN_4; // @[TensorStore.scala 89:23:@24294.6]
  wire  _T_742; // @[Conditional.scala 37:30:@24314.6]
  wire [2:0] _GEN_5; // @[TensorStore.scala 101:33:@24316.8]
  wire  _T_743; // @[Conditional.scala 37:30:@24321.8]
  wire  _T_744; // @[TensorStore.scala 107:19:@24324.12]
  wire  _T_746; // @[TensorStore.scala 109:24:@24329.14]
  wire [2:0] _GEN_6; // @[TensorStore.scala 109:49:@24330.14]
  wire [2:0] _GEN_7; // @[TensorStore.scala 107:29:@24325.12]
  wire [2:0] _GEN_8; // @[TensorStore.scala 106:34:@24323.10]
  wire  _T_747; // @[Conditional.scala 37:30:@24336.10]
  wire  _T_748; // @[Conditional.scala 37:30:@24341.12]
  wire  _T_750; // @[TensorStore.scala 119:19:@24344.16]
  wire [16:0] _T_752; // @[TensorStore.scala 120:31:@24346.18]
  wire [16:0] _T_753; // @[TensorStore.scala 120:31:@24347.18]
  wire [15:0] _T_754; // @[TensorStore.scala 120:31:@24348.18]
  wire  _T_755; // @[TensorStore.scala 120:21:@24349.18]
  wire [16:0] _GEN_103; // @[TensorStore.scala 125:24:@24356.20]
  wire  _T_756; // @[TensorStore.scala 125:24:@24356.20]
  wire [9:0] _T_759; // @[TensorStore.scala 129:42:@24362.22]
  wire [9:0] _T_760; // @[TensorStore.scala 129:42:@24363.22]
  wire [8:0] _T_761; // @[TensorStore.scala 129:42:@24364.22]
  wire [17:0] _T_762; // @[TensorStore.scala 130:29:@24366.22]
  wire [17:0] _T_763; // @[TensorStore.scala 130:29:@24367.22]
  wire [16:0] _T_764; // @[TensorStore.scala 130:29:@24368.22]
  wire [16:0] _GEN_9; // @[TensorStore.scala 125:46:@24357.20]
  wire [16:0] _GEN_10; // @[TensorStore.scala 125:46:@24357.20]
  wire [2:0] _GEN_11; // @[TensorStore.scala 120:38:@24350.18]
  wire [31:0] _GEN_12; // @[TensorStore.scala 120:38:@24350.18]
  wire [16:0] _GEN_13; // @[TensorStore.scala 120:38:@24350.18]
  wire [16:0] _GEN_14; // @[TensorStore.scala 120:38:@24350.18]
  wire [15:0] _GEN_105; // @[TensorStore.scala 134:24:@24374.18]
  wire  _T_765; // @[TensorStore.scala 134:24:@24374.18]
  wire [9:0] _T_768; // @[TensorStore.scala 143:37:@24384.20]
  wire [9:0] _T_769; // @[TensorStore.scala 143:37:@24385.20]
  wire [8:0] _T_770; // @[TensorStore.scala 143:37:@24386.20]
  wire [16:0] _T_771; // @[TensorStore.scala 144:24:@24388.20]
  wire [16:0] _T_772; // @[TensorStore.scala 144:24:@24389.20]
  wire [15:0] _T_773; // @[TensorStore.scala 144:24:@24390.20]
  wire [15:0] _GEN_17; // @[TensorStore.scala 134:45:@24375.18]
  wire [15:0] _GEN_18; // @[TensorStore.scala 134:45:@24375.18]
  wire [2:0] _GEN_19; // @[TensorStore.scala 119:28:@24345.16]
  wire [31:0] _GEN_20; // @[TensorStore.scala 119:28:@24345.16]
  wire [16:0] _GEN_21; // @[TensorStore.scala 119:28:@24345.16]
  wire [16:0] _GEN_22; // @[TensorStore.scala 119:28:@24345.16]
  wire [2:0] _GEN_23; // @[TensorStore.scala 118:27:@24343.14]
  wire [31:0] _GEN_24; // @[TensorStore.scala 118:27:@24343.14]
  wire [16:0] _GEN_25; // @[TensorStore.scala 118:27:@24343.14]
  wire [16:0] _GEN_26; // @[TensorStore.scala 118:27:@24343.14]
  wire [2:0] _GEN_27; // @[Conditional.scala 39:67:@24342.12]
  wire [31:0] _GEN_28; // @[Conditional.scala 39:67:@24342.12]
  wire [16:0] _GEN_29; // @[Conditional.scala 39:67:@24342.12]
  wire [16:0] _GEN_30; // @[Conditional.scala 39:67:@24342.12]
  wire [2:0] _GEN_31; // @[Conditional.scala 39:67:@24337.10]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67:@24337.10]
  wire [16:0] _GEN_33; // @[Conditional.scala 39:67:@24337.10]
  wire [16:0] _GEN_34; // @[Conditional.scala 39:67:@24337.10]
  wire [2:0] _GEN_35; // @[Conditional.scala 39:67:@24322.8]
  wire [31:0] _GEN_36; // @[Conditional.scala 39:67:@24322.8]
  wire [16:0] _GEN_37; // @[Conditional.scala 39:67:@24322.8]
  wire [16:0] _GEN_38; // @[Conditional.scala 39:67:@24322.8]
  wire [2:0] _GEN_39; // @[Conditional.scala 39:67:@24315.6]
  wire [31:0] _GEN_40; // @[Conditional.scala 39:67:@24315.6]
  wire [16:0] _GEN_41; // @[Conditional.scala 39:67:@24315.6]
  wire [16:0] _GEN_42; // @[Conditional.scala 39:67:@24315.6]
  wire [2:0] _GEN_44; // @[Conditional.scala 40:58:@24292.4]
  wire [16:0] _GEN_45; // @[Conditional.scala 40:58:@24292.4]
  wire [16:0] _GEN_46; // @[Conditional.scala 40:58:@24292.4]
  wire [63:0] _T_804; // @[TensorStore.scala 163:46:@24408.4]
  wire [127:0] _T_812; // @[TensorStore.scala 163:46:@24416.4]
  wire  _T_844; // @[TensorStore.scala 170:22:@24433.4]
  wire  _T_845; // @[TensorStore.scala 170:36:@24434.4]
  wire [8:0] _T_847; // @[TensorStore.scala 172:19:@24435.4]
  wire [7:0] _T_848; // @[TensorStore.scala 172:19:@24436.4]
  wire  _T_849; // @[TensorStore.scala 172:10:@24437.4]
  wire  _T_850; // @[TensorStore.scala 171:19:@24438.4]
  wire  _T_853; // @[TensorStore.scala 172:25:@24440.4]
  wire  _T_858; // @[TensorStore.scala 174:10:@24444.4]
  wire  stride; // @[TensorStore.scala 173:18:@24445.4]
  wire  _T_859; // @[TensorStore.scala 176:14:@24446.4]
  wire [16:0] _T_862; // @[TensorStore.scala 179:18:@24452.8]
  wire [15:0] _T_863; // @[TensorStore.scala 179:18:@24453.8]
  wire [15:0] _GEN_58; // @[TensorStore.scala 178:22:@24451.6]
  wire  _T_864; // @[TensorStore.scala 182:14:@24456.4]
  wire  _T_867; // @[TensorStore.scala 182:28:@24458.4]
  wire  _T_869; // @[Decoupled.scala 37:37:@24463.6]
  wire [8:0] _T_871; // @[TensorStore.scala 185:16:@24465.8]
  wire [7:0] _T_872; // @[TensorStore.scala 185:16:@24466.8]
  wire [7:0] _GEN_60; // @[TensorStore.scala 184:37:@24464.6]
  wire  _T_875; // @[TensorStore.scala 189:33:@24470.4]
  wire  _T_878; // @[TensorStore.scala 189:58:@24472.4]
  wire  _T_879; // @[TensorStore.scala 189:25:@24473.4]
  wire  _T_884; // @[TensorStore.scala 191:36:@24480.6]
  wire [8:0] _T_886; // @[TensorStore.scala 192:16:@24482.8]
  wire [7:0] _T_887; // @[TensorStore.scala 192:16:@24483.8]
  wire [7:0] _GEN_62; // @[TensorStore.scala 191:68:@24481.6]
  reg [10:0] raddr_cur; // @[TensorStore.scala 195:22:@24486.4]
  reg [31:0] _RAND_12;
  reg [10:0] raddr_nxt; // @[TensorStore.scala 196:22:@24487.4]
  reg [31:0] _RAND_13;
  wire  _T_894; // @[TensorStore.scala 200:36:@24496.6]
  wire  _T_897; // @[TensorStore.scala 200:68:@24498.6]
  wire [11:0] _T_899; // @[TensorStore.scala 201:28:@24500.8]
  wire [10:0] _T_900; // @[TensorStore.scala 201:28:@24501.8]
  wire [15:0] _GEN_107; // @[TensorStore.scala 203:28:@24506.10]
  wire [16:0] _T_901; // @[TensorStore.scala 203:28:@24506.10]
  wire [15:0] _T_902; // @[TensorStore.scala 203:28:@24507.10]
  wire [15:0] _GEN_64; // @[TensorStore.scala 202:22:@24505.8]
  wire [15:0] _GEN_65; // @[TensorStore.scala 202:22:@24505.8]
  wire [15:0] _GEN_66; // @[TensorStore.scala 200:100:@24499.6]
  wire [15:0] _GEN_67; // @[TensorStore.scala 200:100:@24499.6]
  wire [15:0] _GEN_68; // @[TensorStore.scala 197:25:@24489.4]
  wire [15:0] _GEN_69; // @[TensorStore.scala 197:25:@24489.4]
  wire  _T_907; // @[TensorStore.scala 209:65:@24514.4]
  wire  _T_908; // @[TensorStore.scala 209:57:@24515.4]
  wire  _GEN_71; // @[TensorStore.scala 209:25:@24518.4]
  wire  _T_960; // @[Mux.scala 46:19:@24531.4]
  wire [63:0] mdata_0; // @[Mux.scala 46:16:@24532.4]
  wire [63:0] mdata_1; // @[Mux.scala 46:16:@24532.4]
  wire  _T_975; // @[TensorStore.scala 217:59:@24541.6]
  wire  _T_976; // @[TensorStore.scala 217:51:@24542.6]
  wire [31:0] _GEN_74; // @[TensorStore.scala 219:22:@24547.8]
  wire [31:0] _GEN_75; // @[TensorStore.scala 219:22:@24547.8]
  wire [31:0] _GEN_76; // @[TensorStore.scala 217:68:@24543.6]
  wire [31:0] _GEN_77; // @[TensorStore.scala 217:68:@24543.6]
  wire [35:0] _GEN_78; // @[TensorStore.scala 214:25:@24534.4]
  wire [35:0] _GEN_79; // @[TensorStore.scala 214:25:@24534.4]
  wire  _T_982; // @[:@24557.4]
  wire [8:0] _T_987; // @[TensorStore.scala 234:18:@24566.8]
  wire [7:0] _T_988; // @[TensorStore.scala 234:18:@24567.8]
  wire [7:0] _GEN_82; // @[TensorStore.scala 233:37:@24565.6]
  wire  _T_1010; // @[TensorStore.scala 241:50:@24590.4]
  reg [10:0] tensorFile_0_0__T_914_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [10:0] tensorFile_0_1__T_914_addr_pipe_0;
  reg [31:0] _RAND_15;
  assign tensorFile_0_0__T_914_addr = tensorFile_0_0__T_914_addr_pipe_0;
  assign tensorFile_0_0__T_914_data = tensorFile_0_0[tensorFile_0_0__T_914_addr]; // @[TensorStore.scala 152:16:@24395.4]
  assign tensorFile_0_0__T_836_data = _T_812[63:0];
  assign tensorFile_0_0__T_836_addr = io_tensor_wr_bits_idx;
  assign tensorFile_0_0__T_836_mask = 1'h1;
  assign tensorFile_0_0__T_836_en = io_tensor_wr_valid;
  assign tensorFile_0_1__T_914_addr = tensorFile_0_1__T_914_addr_pipe_0;
  assign tensorFile_0_1__T_914_data = tensorFile_0_1[tensorFile_0_1__T_914_addr]; // @[TensorStore.scala 152:16:@24395.4]
  assign tensorFile_0_1__T_836_data = _T_812[127:64];
  assign tensorFile_0_1__T_836_addr = io_tensor_wr_bits_idx;
  assign tensorFile_0_1__T_836_mask = 1'h1;
  assign tensorFile_0_1__T_836_en = io_tensor_wr_valid;
  assign dec_sram_offset = io_inst[24:9]; // @[TensorStore.scala 51:29:@24170.4]
  assign dec_dram_offset = io_inst[56:25]; // @[TensorStore.scala 51:29:@24172.4]
  assign dec_ysize = io_inst[79:64]; // @[TensorStore.scala 51:29:@24176.4]
  assign dec_xsize = io_inst[95:80]; // @[TensorStore.scala 51:29:@24178.4]
  assign dec_xstride = io_inst[111:96]; // @[TensorStore.scala 51:29:@24180.4]
  assign _GEN_96 = {{1'd0}, dec_xsize}; // @[TensorStore.scala 57:26:@24195.4]
  assign _T_610 = _GEN_96 << 1; // @[TensorStore.scala 57:26:@24195.4]
  assign _T_612 = _T_610 - 17'h1; // @[TensorStore.scala 57:67:@24196.4]
  assign _T_613 = $unsigned(_T_612); // @[TensorStore.scala 57:67:@24197.4]
  assign xsize = _T_613[16:0]; // @[TensorStore.scala 57:67:@24198.4]
  assign _GEN_97 = {{4'd0}, dec_xstride}; // @[TensorStore.scala 66:35:@24203.4]
  assign xstride_bytes = _GEN_97 << 4; // @[TensorStore.scala 66:35:@24203.4]
  assign _GEN_98 = {{4'd0}, dec_dram_offset}; // @[TensorStore.scala 71:66:@24268.4]
  assign _T_718 = _GEN_98 << 4; // @[TensorStore.scala 71:66:@24268.4]
  assign _T_719 = 36'hffffffff & _T_718; // @[TensorStore.scala 71:47:@24269.4]
  assign _GEN_99 = {{4'd0}, io_baddr}; // @[TensorStore.scala 71:33:@24270.4]
  assign xfer_init_addr = _GEN_99 | _T_719; // @[TensorStore.scala 71:33:@24270.4]
  assign _T_720 = waddr_cur + xfer_bytes; // @[TensorStore.scala 72:35:@24271.4]
  assign xfer_split_addr = waddr_cur + xfer_bytes; // @[TensorStore.scala 72:35:@24272.4]
  assign _GEN_100 = {{12'd0}, xstride_bytes}; // @[TensorStore.scala 73:36:@24273.4]
  assign _T_721 = waddr_nxt + _GEN_100; // @[TensorStore.scala 73:36:@24273.4]
  assign xfer_stride_addr = waddr_nxt + _GEN_100; // @[TensorStore.scala 73:36:@24274.4]
  assign _GEN_15 = xfer_init_addr % 36'h800; // @[TensorStore.scala 75:55:@24275.4]
  assign _T_722 = _GEN_15[11:0]; // @[TensorStore.scala 75:55:@24275.4]
  assign _T_723 = 12'h800 - _T_722; // @[TensorStore.scala 75:38:@24276.4]
  assign _T_724 = $unsigned(_T_723); // @[TensorStore.scala 75:38:@24277.4]
  assign xfer_init_bytes = _T_724[11:0]; // @[TensorStore.scala 75:38:@24278.4]
  assign xfer_init_pulses = xfer_init_bytes[11:3]; // @[TensorStore.scala 76:43:@24279.4]
  assign _GEN_16 = xfer_split_addr % 32'h800; // @[TensorStore.scala 77:56:@24280.4]
  assign _T_725 = _GEN_16[11:0]; // @[TensorStore.scala 77:56:@24280.4]
  assign _T_726 = 12'h800 - _T_725; // @[TensorStore.scala 77:38:@24281.4]
  assign _T_727 = $unsigned(_T_726); // @[TensorStore.scala 77:38:@24282.4]
  assign xfer_split_bytes = _T_727[11:0]; // @[TensorStore.scala 77:38:@24283.4]
  assign xfer_split_pulses = xfer_split_bytes[11:3]; // @[TensorStore.scala 78:44:@24284.4]
  assign _GEN_43 = xfer_stride_addr % 32'h800; // @[TensorStore.scala 79:57:@24285.4]
  assign _T_728 = _GEN_43[11:0]; // @[TensorStore.scala 79:57:@24285.4]
  assign _T_729 = 12'h800 - _T_728; // @[TensorStore.scala 79:38:@24286.4]
  assign _T_730 = $unsigned(_T_729); // @[TensorStore.scala 79:38:@24287.4]
  assign xfer_stride_bytes = _T_730[11:0]; // @[TensorStore.scala 79:38:@24288.4]
  assign xfer_stride_pulses = xfer_stride_bytes[11:3]; // @[TensorStore.scala 80:45:@24289.4]
  assign _T_732 = 3'h0 == state; // @[Conditional.scala 37:30:@24291.4]
  assign _GEN_101 = {{8'd0}, xfer_init_pulses}; // @[TensorStore.scala 91:21:@24296.8]
  assign _T_733 = xsize < _GEN_101; // @[TensorStore.scala 91:21:@24296.8]
  assign _T_736 = xfer_init_pulses - 9'h1; // @[TensorStore.scala 95:36:@24302.10]
  assign _T_737 = $unsigned(_T_736); // @[TensorStore.scala 95:36:@24303.10]
  assign _T_738 = _T_737[8:0]; // @[TensorStore.scala 95:36:@24304.10]
  assign _T_739 = xsize - _GEN_101; // @[TensorStore.scala 96:25:@24306.10]
  assign _T_740 = $unsigned(_T_739); // @[TensorStore.scala 96:25:@24307.10]
  assign _T_741 = _T_740[16:0]; // @[TensorStore.scala 96:25:@24308.10]
  assign _GEN_0 = _T_733 ? xsize : {{8'd0}, _T_738}; // @[TensorStore.scala 91:41:@24297.8]
  assign _GEN_1 = _T_733 ? 17'h0 : _T_741; // @[TensorStore.scala 91:41:@24297.8]
  assign _GEN_2 = io_start ? 3'h1 : state; // @[TensorStore.scala 89:23:@24294.6]
  assign _GEN_3 = io_start ? _GEN_0 : {{9'd0}, xlen}; // @[TensorStore.scala 89:23:@24294.6]
  assign _GEN_4 = io_start ? _GEN_1 : {{1'd0}, xrem}; // @[TensorStore.scala 89:23:@24294.6]
  assign _T_742 = 3'h1 == state; // @[Conditional.scala 37:30:@24314.6]
  assign _GEN_5 = io_vme_wr_cmd_ready ? 3'h2 : state; // @[TensorStore.scala 101:33:@24316.8]
  assign _T_743 = 3'h2 == state; // @[Conditional.scala 37:30:@24321.8]
  assign _T_744 = xcnt == xlen; // @[TensorStore.scala 107:19:@24324.12]
  assign _T_746 = tag == 8'h1; // @[TensorStore.scala 109:24:@24329.14]
  assign _GEN_6 = _T_746 ? 3'h3 : state; // @[TensorStore.scala 109:49:@24330.14]
  assign _GEN_7 = _T_744 ? 3'h4 : _GEN_6; // @[TensorStore.scala 107:29:@24325.12]
  assign _GEN_8 = io_vme_wr_data_ready ? _GEN_7 : state; // @[TensorStore.scala 106:34:@24323.10]
  assign _T_747 = 3'h3 == state; // @[Conditional.scala 37:30:@24336.10]
  assign _T_748 = 3'h4 == state; // @[Conditional.scala 37:30:@24341.12]
  assign _T_750 = xrem == 16'h0; // @[TensorStore.scala 119:19:@24344.16]
  assign _T_752 = dec_ysize - 16'h1; // @[TensorStore.scala 120:31:@24346.18]
  assign _T_753 = $unsigned(_T_752); // @[TensorStore.scala 120:31:@24347.18]
  assign _T_754 = _T_753[15:0]; // @[TensorStore.scala 120:31:@24348.18]
  assign _T_755 = ycnt == _T_754; // @[TensorStore.scala 120:21:@24349.18]
  assign _GEN_103 = {{8'd0}, xfer_stride_pulses}; // @[TensorStore.scala 125:24:@24356.20]
  assign _T_756 = xsize < _GEN_103; // @[TensorStore.scala 125:24:@24356.20]
  assign _T_759 = xfer_stride_pulses - 9'h1; // @[TensorStore.scala 129:42:@24362.22]
  assign _T_760 = $unsigned(_T_759); // @[TensorStore.scala 129:42:@24363.22]
  assign _T_761 = _T_760[8:0]; // @[TensorStore.scala 129:42:@24364.22]
  assign _T_762 = xsize - _GEN_103; // @[TensorStore.scala 130:29:@24366.22]
  assign _T_763 = $unsigned(_T_762); // @[TensorStore.scala 130:29:@24367.22]
  assign _T_764 = _T_763[16:0]; // @[TensorStore.scala 130:29:@24368.22]
  assign _GEN_9 = _T_756 ? xsize : {{8'd0}, _T_761}; // @[TensorStore.scala 125:46:@24357.20]
  assign _GEN_10 = _T_756 ? 17'h0 : _T_764; // @[TensorStore.scala 125:46:@24357.20]
  assign _GEN_11 = _T_755 ? 3'h0 : 3'h1; // @[TensorStore.scala 120:38:@24350.18]
  assign _GEN_12 = _T_755 ? xfer_bytes : {{20'd0}, xfer_stride_bytes}; // @[TensorStore.scala 120:38:@24350.18]
  assign _GEN_13 = _T_755 ? {{9'd0}, xlen} : _GEN_9; // @[TensorStore.scala 120:38:@24350.18]
  assign _GEN_14 = _T_755 ? {{1'd0}, xrem} : _GEN_10; // @[TensorStore.scala 120:38:@24350.18]
  assign _GEN_105 = {{7'd0}, xfer_split_pulses}; // @[TensorStore.scala 134:24:@24374.18]
  assign _T_765 = xrem < _GEN_105; // @[TensorStore.scala 134:24:@24374.18]
  assign _T_768 = xfer_split_pulses - 9'h1; // @[TensorStore.scala 143:37:@24384.20]
  assign _T_769 = $unsigned(_T_768); // @[TensorStore.scala 143:37:@24385.20]
  assign _T_770 = _T_769[8:0]; // @[TensorStore.scala 143:37:@24386.20]
  assign _T_771 = xrem - _GEN_105; // @[TensorStore.scala 144:24:@24388.20]
  assign _T_772 = $unsigned(_T_771); // @[TensorStore.scala 144:24:@24389.20]
  assign _T_773 = _T_772[15:0]; // @[TensorStore.scala 144:24:@24390.20]
  assign _GEN_17 = _T_765 ? xrem : {{7'd0}, _T_770}; // @[TensorStore.scala 134:45:@24375.18]
  assign _GEN_18 = _T_765 ? 16'h0 : _T_773; // @[TensorStore.scala 134:45:@24375.18]
  assign _GEN_19 = _T_750 ? _GEN_11 : 3'h1; // @[TensorStore.scala 119:28:@24345.16]
  assign _GEN_20 = _T_750 ? _GEN_12 : {{20'd0}, xfer_split_bytes}; // @[TensorStore.scala 119:28:@24345.16]
  assign _GEN_21 = _T_750 ? _GEN_13 : {{1'd0}, _GEN_17}; // @[TensorStore.scala 119:28:@24345.16]
  assign _GEN_22 = _T_750 ? _GEN_14 : {{1'd0}, _GEN_18}; // @[TensorStore.scala 119:28:@24345.16]
  assign _GEN_23 = io_vme_wr_ack ? _GEN_19 : state; // @[TensorStore.scala 118:27:@24343.14]
  assign _GEN_24 = io_vme_wr_ack ? _GEN_20 : xfer_bytes; // @[TensorStore.scala 118:27:@24343.14]
  assign _GEN_25 = io_vme_wr_ack ? _GEN_21 : {{9'd0}, xlen}; // @[TensorStore.scala 118:27:@24343.14]
  assign _GEN_26 = io_vme_wr_ack ? _GEN_22 : {{1'd0}, xrem}; // @[TensorStore.scala 118:27:@24343.14]
  assign _GEN_27 = _T_748 ? _GEN_23 : state; // @[Conditional.scala 39:67:@24342.12]
  assign _GEN_28 = _T_748 ? _GEN_24 : xfer_bytes; // @[Conditional.scala 39:67:@24342.12]
  assign _GEN_29 = _T_748 ? _GEN_25 : {{9'd0}, xlen}; // @[Conditional.scala 39:67:@24342.12]
  assign _GEN_30 = _T_748 ? _GEN_26 : {{1'd0}, xrem}; // @[Conditional.scala 39:67:@24342.12]
  assign _GEN_31 = _T_747 ? 3'h2 : _GEN_27; // @[Conditional.scala 39:67:@24337.10]
  assign _GEN_32 = _T_747 ? xfer_bytes : _GEN_28; // @[Conditional.scala 39:67:@24337.10]
  assign _GEN_33 = _T_747 ? {{9'd0}, xlen} : _GEN_29; // @[Conditional.scala 39:67:@24337.10]
  assign _GEN_34 = _T_747 ? {{1'd0}, xrem} : _GEN_30; // @[Conditional.scala 39:67:@24337.10]
  assign _GEN_35 = _T_743 ? _GEN_8 : _GEN_31; // @[Conditional.scala 39:67:@24322.8]
  assign _GEN_36 = _T_743 ? xfer_bytes : _GEN_32; // @[Conditional.scala 39:67:@24322.8]
  assign _GEN_37 = _T_743 ? {{9'd0}, xlen} : _GEN_33; // @[Conditional.scala 39:67:@24322.8]
  assign _GEN_38 = _T_743 ? {{1'd0}, xrem} : _GEN_34; // @[Conditional.scala 39:67:@24322.8]
  assign _GEN_39 = _T_742 ? _GEN_5 : _GEN_35; // @[Conditional.scala 39:67:@24315.6]
  assign _GEN_40 = _T_742 ? xfer_bytes : _GEN_36; // @[Conditional.scala 39:67:@24315.6]
  assign _GEN_41 = _T_742 ? {{9'd0}, xlen} : _GEN_37; // @[Conditional.scala 39:67:@24315.6]
  assign _GEN_42 = _T_742 ? {{1'd0}, xrem} : _GEN_38; // @[Conditional.scala 39:67:@24315.6]
  assign _GEN_44 = _T_732 ? _GEN_2 : _GEN_39; // @[Conditional.scala 40:58:@24292.4]
  assign _GEN_45 = _T_732 ? _GEN_3 : _GEN_41; // @[Conditional.scala 40:58:@24292.4]
  assign _GEN_46 = _T_732 ? _GEN_4 : _GEN_42; // @[Conditional.scala 40:58:@24292.4]
  assign _T_804 = {io_tensor_wr_bits_data_0_7,io_tensor_wr_bits_data_0_6,io_tensor_wr_bits_data_0_5,io_tensor_wr_bits_data_0_4,io_tensor_wr_bits_data_0_3,io_tensor_wr_bits_data_0_2,io_tensor_wr_bits_data_0_1,io_tensor_wr_bits_data_0_0}; // @[TensorStore.scala 163:46:@24408.4]
  assign _T_812 = {io_tensor_wr_bits_data_0_15,io_tensor_wr_bits_data_0_14,io_tensor_wr_bits_data_0_13,io_tensor_wr_bits_data_0_12,io_tensor_wr_bits_data_0_11,io_tensor_wr_bits_data_0_10,io_tensor_wr_bits_data_0_9,io_tensor_wr_bits_data_0_8,_T_804}; // @[TensorStore.scala 163:46:@24416.4]
  assign _T_844 = state == 3'h4; // @[TensorStore.scala 170:22:@24433.4]
  assign _T_845 = _T_844 & io_vme_wr_ack; // @[TensorStore.scala 170:36:@24434.4]
  assign _T_847 = xlen + 8'h1; // @[TensorStore.scala 172:19:@24435.4]
  assign _T_848 = xlen + 8'h1; // @[TensorStore.scala 172:19:@24436.4]
  assign _T_849 = xcnt == _T_848; // @[TensorStore.scala 172:10:@24437.4]
  assign _T_850 = _T_845 & _T_849; // @[TensorStore.scala 171:19:@24438.4]
  assign _T_853 = _T_850 & _T_750; // @[TensorStore.scala 172:25:@24440.4]
  assign _T_858 = ycnt != _T_754; // @[TensorStore.scala 174:10:@24444.4]
  assign stride = _T_853 & _T_858; // @[TensorStore.scala 173:18:@24445.4]
  assign _T_859 = state == 3'h0; // @[TensorStore.scala 176:14:@24446.4]
  assign _T_862 = ycnt + 16'h1; // @[TensorStore.scala 179:18:@24452.8]
  assign _T_863 = ycnt + 16'h1; // @[TensorStore.scala 179:18:@24453.8]
  assign _GEN_58 = stride ? _T_863 : ycnt; // @[TensorStore.scala 178:22:@24451.6]
  assign _T_864 = state == 3'h1; // @[TensorStore.scala 182:14:@24456.4]
  assign _T_867 = _T_864 | _T_746; // @[TensorStore.scala 182:28:@24458.4]
  assign _T_869 = io_vme_wr_data_ready & io_vme_wr_data_valid; // @[Decoupled.scala 37:37:@24463.6]
  assign _T_871 = tag + 8'h1; // @[TensorStore.scala 185:16:@24465.8]
  assign _T_872 = tag + 8'h1; // @[TensorStore.scala 185:16:@24466.8]
  assign _GEN_60 = _T_869 ? _T_872 : tag; // @[TensorStore.scala 184:37:@24464.6]
  assign _T_875 = set == 8'h0; // @[TensorStore.scala 189:33:@24470.4]
  assign _T_878 = _T_875 & _T_746; // @[TensorStore.scala 189:58:@24472.4]
  assign _T_879 = _T_864 | _T_878; // @[TensorStore.scala 189:25:@24473.4]
  assign _T_884 = _T_869 & _T_746; // @[TensorStore.scala 191:36:@24480.6]
  assign _T_886 = set + 8'h1; // @[TensorStore.scala 192:16:@24482.8]
  assign _T_887 = set + 8'h1; // @[TensorStore.scala 192:16:@24483.8]
  assign _GEN_62 = _T_884 ? _T_887 : set; // @[TensorStore.scala 191:68:@24481.6]
  assign _T_894 = _T_869 & _T_875; // @[TensorStore.scala 200:36:@24496.6]
  assign _T_897 = _T_894 & _T_746; // @[TensorStore.scala 200:68:@24498.6]
  assign _T_899 = raddr_cur + 11'h1; // @[TensorStore.scala 201:28:@24500.8]
  assign _T_900 = raddr_cur + 11'h1; // @[TensorStore.scala 201:28:@24501.8]
  assign _GEN_107 = {{5'd0}, raddr_nxt}; // @[TensorStore.scala 203:28:@24506.10]
  assign _T_901 = _GEN_107 + dec_xsize; // @[TensorStore.scala 203:28:@24506.10]
  assign _T_902 = _GEN_107 + dec_xsize; // @[TensorStore.scala 203:28:@24507.10]
  assign _GEN_64 = stride ? _T_902 : {{5'd0}, raddr_cur}; // @[TensorStore.scala 202:22:@24505.8]
  assign _GEN_65 = stride ? _T_902 : {{5'd0}, raddr_nxt}; // @[TensorStore.scala 202:22:@24505.8]
  assign _GEN_66 = _T_897 ? {{5'd0}, _T_900} : _GEN_64; // @[TensorStore.scala 200:100:@24499.6]
  assign _GEN_67 = _T_897 ? {{5'd0}, raddr_nxt} : _GEN_65; // @[TensorStore.scala 200:100:@24499.6]
  assign _GEN_68 = _T_859 ? dec_sram_offset : _GEN_66; // @[TensorStore.scala 197:25:@24489.4]
  assign _GEN_69 = _T_859 ? dec_sram_offset : _GEN_67; // @[TensorStore.scala 197:25:@24489.4]
  assign _T_907 = state == 3'h3; // @[TensorStore.scala 209:65:@24514.4]
  assign _T_908 = _T_864 | _T_907; // @[TensorStore.scala 209:57:@24515.4]
  assign _GEN_71 = _T_908; // @[TensorStore.scala 209:25:@24518.4]
  assign _T_960 = 8'h0 == set; // @[Mux.scala 46:19:@24531.4]
  assign mdata_0 = _T_960 ? tensorFile_0_0__T_914_data : 64'h0; // @[Mux.scala 46:16:@24532.4]
  assign mdata_1 = _T_960 ? tensorFile_0_1__T_914_data : 64'h0; // @[Mux.scala 46:16:@24532.4]
  assign _T_975 = xrem != 16'h0; // @[TensorStore.scala 217:59:@24541.6]
  assign _T_976 = _T_845 & _T_975; // @[TensorStore.scala 217:51:@24542.6]
  assign _GEN_74 = stride ? xfer_stride_addr : waddr_cur; // @[TensorStore.scala 219:22:@24547.8]
  assign _GEN_75 = stride ? xfer_stride_addr : waddr_nxt; // @[TensorStore.scala 219:22:@24547.8]
  assign _GEN_76 = _T_976 ? xfer_split_addr : _GEN_74; // @[TensorStore.scala 217:68:@24543.6]
  assign _GEN_77 = _T_976 ? waddr_nxt : _GEN_75; // @[TensorStore.scala 217:68:@24543.6]
  assign _GEN_78 = _T_859 ? xfer_init_addr : {{4'd0}, _GEN_76}; // @[TensorStore.scala 214:25:@24534.4]
  assign _GEN_79 = _T_859 ? xfer_init_addr : {{4'd0}, _GEN_77}; // @[TensorStore.scala 214:25:@24534.4]
  assign _T_982 = tag[0]; // @[:@24557.4]
  assign _T_987 = xcnt + 8'h1; // @[TensorStore.scala 234:18:@24566.8]
  assign _T_988 = xcnt + 8'h1; // @[TensorStore.scala 234:18:@24567.8]
  assign _GEN_82 = _T_869 ? _T_988 : xcnt; // @[TensorStore.scala 233:37:@24565.6]
  assign _T_1010 = _T_845 & _T_750; // @[TensorStore.scala 241:50:@24590.4]
  assign io_done = _T_1010 & _T_755; // @[TensorStore.scala 241:11:@24596.4]
  assign io_vme_wr_cmd_valid = state == 3'h1; // @[TensorStore.scala 224:23:@24552.4]
  assign io_vme_wr_cmd_bits_addr = waddr_cur; // @[TensorStore.scala 225:27:@24553.4]
  assign io_vme_wr_cmd_bits_len = xlen; // @[TensorStore.scala 226:26:@24554.4]
  assign io_vme_wr_data_valid = state == 3'h2; // @[TensorStore.scala 228:24:@24556.4]
  assign io_vme_wr_data_bits = _T_982 ? mdata_1 : mdata_0; // @[TensorStore.scala 229:23:@24558.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_0[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    tensorFile_0_1[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  waddr_cur = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  waddr_nxt = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  xcnt = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  xlen = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  xrem = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ycnt = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tag = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  set = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  xfer_bytes = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  raddr_cur = _RAND_12[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  raddr_nxt = _RAND_13[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  tensorFile_0_0__T_914_addr_pipe_0 = _RAND_14[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  tensorFile_0_1__T_914_addr_pipe_0 = _RAND_15[10:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tensorFile_0_0__T_836_en & tensorFile_0_0__T_836_mask) begin
      tensorFile_0_0[tensorFile_0_0__T_836_addr] <= tensorFile_0_0__T_836_data; // @[TensorStore.scala 152:16:@24395.4]
    end
    if(tensorFile_0_1__T_836_en & tensorFile_0_1__T_836_mask) begin
      tensorFile_0_1[tensorFile_0_1__T_836_addr] <= tensorFile_0_1__T_836_data; // @[TensorStore.scala 152:16:@24395.4]
    end
    waddr_cur <= _GEN_78[31:0];
    waddr_nxt <= _GEN_79[31:0];
    if (_T_864) begin
      xcnt <= 8'h0;
    end else begin
      if (_T_869) begin
        xcnt <= _T_988;
      end
    end
    xlen <= _GEN_45[7:0];
    xrem <= _GEN_46[15:0];
    if (_T_859) begin
      ycnt <= 16'h0;
    end else begin
      if (stride) begin
        ycnt <= _T_863;
      end
    end
    if (_T_867) begin
      tag <= 8'h0;
    end else begin
      if (_T_869) begin
        tag <= _T_872;
      end
    end
    if (_T_879) begin
      set <= 8'h0;
    end else begin
      if (_T_884) begin
        set <= _T_887;
      end
    end
    if (_T_732) begin
      xfer_bytes <= {{20'd0}, xfer_init_bytes};
    end else begin
      if (!(_T_742)) begin
        if (!(_T_743)) begin
          if (!(_T_747)) begin
            if (_T_748) begin
              if (io_vme_wr_ack) begin
                if (_T_750) begin
                  if (!(_T_755)) begin
                    xfer_bytes <= {{20'd0}, xfer_stride_bytes};
                  end
                end else begin
                  xfer_bytes <= {{20'd0}, xfer_split_bytes};
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_732) begin
        if (io_start) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_742) begin
          if (io_vme_wr_cmd_ready) begin
            state <= 3'h2;
          end
        end else begin
          if (_T_743) begin
            if (io_vme_wr_data_ready) begin
              if (_T_744) begin
                state <= 3'h4;
              end else begin
                if (_T_746) begin
                  state <= 3'h3;
                end
              end
            end
          end else begin
            if (_T_747) begin
              state <= 3'h2;
            end else begin
              if (_T_748) begin
                if (io_vme_wr_ack) begin
                  if (_T_750) begin
                    if (_T_755) begin
                      state <= 3'h0;
                    end else begin
                      state <= 3'h1;
                    end
                  end else begin
                    state <= 3'h1;
                  end
                end
              end
            end
          end
        end
      end
    end
    raddr_cur <= _GEN_68[10:0];
    raddr_nxt <= _GEN_69[10:0];
    if (_GEN_71) begin
      tensorFile_0_0__T_914_addr_pipe_0 <= raddr_cur;
    end
    if (_GEN_71) begin
      tensorFile_0_1__T_914_addr_pipe_0 <= raddr_cur;
    end
  end
endmodule
module Store( // @[:@24598.2]
  input          clock, // @[:@24599.4]
  input          reset, // @[:@24600.4]
  input          io_i_post, // @[:@24601.4]
  output         io_o_post, // @[:@24601.4]
  output         io_inst_ready, // @[:@24601.4]
  input          io_inst_valid, // @[:@24601.4]
  input  [127:0] io_inst_bits, // @[:@24601.4]
  input  [31:0]  io_out_baddr, // @[:@24601.4]
  input          io_vme_wr_cmd_ready, // @[:@24601.4]
  output         io_vme_wr_cmd_valid, // @[:@24601.4]
  output [31:0]  io_vme_wr_cmd_bits_addr, // @[:@24601.4]
  output [7:0]   io_vme_wr_cmd_bits_len, // @[:@24601.4]
  input          io_vme_wr_data_ready, // @[:@24601.4]
  output         io_vme_wr_data_valid, // @[:@24601.4]
  output [63:0]  io_vme_wr_data_bits, // @[:@24601.4]
  input          io_vme_wr_ack, // @[:@24601.4]
  input          io_out_wr_valid, // @[:@24601.4]
  input  [10:0]  io_out_wr_bits_idx, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_0, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_1, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_2, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_3, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_4, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_5, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_6, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_7, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_8, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_9, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_10, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_11, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_12, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_13, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_14, // @[:@24601.4]
  input  [7:0]   io_out_wr_bits_data_0_15 // @[:@24601.4]
);
  wire  s_clock; // @[Store.scala 46:17:@24604.4]
  wire  s_reset; // @[Store.scala 46:17:@24604.4]
  wire  s_io_spost; // @[Store.scala 46:17:@24604.4]
  wire  s_io_swait; // @[Store.scala 46:17:@24604.4]
  wire  s_io_sready; // @[Store.scala 46:17:@24604.4]
  wire  inst_q_clock; // @[Store.scala 47:22:@24607.4]
  wire  inst_q_reset; // @[Store.scala 47:22:@24607.4]
  wire  inst_q_io_enq_ready; // @[Store.scala 47:22:@24607.4]
  wire  inst_q_io_enq_valid; // @[Store.scala 47:22:@24607.4]
  wire [127:0] inst_q_io_enq_bits; // @[Store.scala 47:22:@24607.4]
  wire  inst_q_io_deq_ready; // @[Store.scala 47:22:@24607.4]
  wire  inst_q_io_deq_valid; // @[Store.scala 47:22:@24607.4]
  wire [127:0] inst_q_io_deq_bits; // @[Store.scala 47:22:@24607.4]
  wire [127:0] dec_io_inst; // @[Store.scala 49:19:@24610.4]
  wire  dec_io_push_prev; // @[Store.scala 49:19:@24610.4]
  wire  dec_io_pop_prev; // @[Store.scala 49:19:@24610.4]
  wire  dec_io_isStore; // @[Store.scala 49:19:@24610.4]
  wire  dec_io_isSync; // @[Store.scala 49:19:@24610.4]
  wire  tensorStore_clock; // @[Store.scala 52:27:@24614.4]
  wire  tensorStore_reset; // @[Store.scala 52:27:@24614.4]
  wire  tensorStore_io_start; // @[Store.scala 52:27:@24614.4]
  wire  tensorStore_io_done; // @[Store.scala 52:27:@24614.4]
  wire [127:0] tensorStore_io_inst; // @[Store.scala 52:27:@24614.4]
  wire [31:0] tensorStore_io_baddr; // @[Store.scala 52:27:@24614.4]
  wire  tensorStore_io_vme_wr_cmd_ready; // @[Store.scala 52:27:@24614.4]
  wire  tensorStore_io_vme_wr_cmd_valid; // @[Store.scala 52:27:@24614.4]
  wire [31:0] tensorStore_io_vme_wr_cmd_bits_addr; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_vme_wr_cmd_bits_len; // @[Store.scala 52:27:@24614.4]
  wire  tensorStore_io_vme_wr_data_ready; // @[Store.scala 52:27:@24614.4]
  wire  tensorStore_io_vme_wr_data_valid; // @[Store.scala 52:27:@24614.4]
  wire [63:0] tensorStore_io_vme_wr_data_bits; // @[Store.scala 52:27:@24614.4]
  wire  tensorStore_io_vme_wr_ack; // @[Store.scala 52:27:@24614.4]
  wire  tensorStore_io_tensor_wr_valid; // @[Store.scala 52:27:@24614.4]
  wire [10:0] tensorStore_io_tensor_wr_bits_idx; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_0; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_1; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_2; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_3; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_4; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_5; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_6; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_7; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_8; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_9; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_10; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_11; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_12; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_13; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_14; // @[Store.scala 52:27:@24614.4]
  wire [7:0] tensorStore_io_tensor_wr_bits_data_0_15; // @[Store.scala 52:27:@24614.4]
  reg [1:0] state; // @[Store.scala 44:22:@24603.4]
  reg [31:0] _RAND_0;
  wire  _T_597; // @[Store.scala 54:40:@24617.4]
  wire  start; // @[Store.scala 54:35:@24618.4]
  wire  _T_598; // @[Conditional.scala 37:30:@24619.4]
  wire [1:0] _GEN_0; // @[Store.scala 63:36:@24626.10]
  wire [1:0] _GEN_1; // @[Store.scala 61:29:@24622.8]
  wire [1:0] _GEN_2; // @[Store.scala 60:19:@24621.6]
  wire  _T_599; // @[Conditional.scala 37:30:@24632.6]
  wire  _T_600; // @[Conditional.scala 37:30:@24637.8]
  wire [1:0] _GEN_3; // @[Store.scala 72:18:@24639.10]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@24638.8]
  wire [1:0] _GEN_5; // @[Conditional.scala 39:67:@24633.6]
  wire [1:0] _GEN_6; // @[Conditional.scala 40:58:@24620.4]
  wire  _T_601; // @[Store.scala 80:33:@24646.4]
  wire  _T_602; // @[Store.scala 80:42:@24647.4]
  wire  _T_603; // @[Store.scala 80:59:@24648.4]
  wire  _T_604; // @[Store.scala 80:50:@24649.4]
  wire  _T_605; // @[Store.scala 83:33:@24651.4]
  wire  _T_606; // @[Store.scala 83:43:@24652.4]
  Semaphore s ( // @[Store.scala 46:17:@24604.4]
    .clock(s_clock),
    .reset(s_reset),
    .io_spost(s_io_spost),
    .io_swait(s_io_swait),
    .io_sready(s_io_sready)
  );
  Queue_1 inst_q ( // @[Store.scala 47:22:@24607.4]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits)
  );
  StoreDecode dec ( // @[Store.scala 49:19:@24610.4]
    .io_inst(dec_io_inst),
    .io_push_prev(dec_io_push_prev),
    .io_pop_prev(dec_io_pop_prev),
    .io_isStore(dec_io_isStore),
    .io_isSync(dec_io_isSync)
  );
  TensorStore tensorStore ( // @[Store.scala 52:27:@24614.4]
    .clock(tensorStore_clock),
    .reset(tensorStore_reset),
    .io_start(tensorStore_io_start),
    .io_done(tensorStore_io_done),
    .io_inst(tensorStore_io_inst),
    .io_baddr(tensorStore_io_baddr),
    .io_vme_wr_cmd_ready(tensorStore_io_vme_wr_cmd_ready),
    .io_vme_wr_cmd_valid(tensorStore_io_vme_wr_cmd_valid),
    .io_vme_wr_cmd_bits_addr(tensorStore_io_vme_wr_cmd_bits_addr),
    .io_vme_wr_cmd_bits_len(tensorStore_io_vme_wr_cmd_bits_len),
    .io_vme_wr_data_ready(tensorStore_io_vme_wr_data_ready),
    .io_vme_wr_data_valid(tensorStore_io_vme_wr_data_valid),
    .io_vme_wr_data_bits(tensorStore_io_vme_wr_data_bits),
    .io_vme_wr_ack(tensorStore_io_vme_wr_ack),
    .io_tensor_wr_valid(tensorStore_io_tensor_wr_valid),
    .io_tensor_wr_bits_idx(tensorStore_io_tensor_wr_bits_idx),
    .io_tensor_wr_bits_data_0_0(tensorStore_io_tensor_wr_bits_data_0_0),
    .io_tensor_wr_bits_data_0_1(tensorStore_io_tensor_wr_bits_data_0_1),
    .io_tensor_wr_bits_data_0_2(tensorStore_io_tensor_wr_bits_data_0_2),
    .io_tensor_wr_bits_data_0_3(tensorStore_io_tensor_wr_bits_data_0_3),
    .io_tensor_wr_bits_data_0_4(tensorStore_io_tensor_wr_bits_data_0_4),
    .io_tensor_wr_bits_data_0_5(tensorStore_io_tensor_wr_bits_data_0_5),
    .io_tensor_wr_bits_data_0_6(tensorStore_io_tensor_wr_bits_data_0_6),
    .io_tensor_wr_bits_data_0_7(tensorStore_io_tensor_wr_bits_data_0_7),
    .io_tensor_wr_bits_data_0_8(tensorStore_io_tensor_wr_bits_data_0_8),
    .io_tensor_wr_bits_data_0_9(tensorStore_io_tensor_wr_bits_data_0_9),
    .io_tensor_wr_bits_data_0_10(tensorStore_io_tensor_wr_bits_data_0_10),
    .io_tensor_wr_bits_data_0_11(tensorStore_io_tensor_wr_bits_data_0_11),
    .io_tensor_wr_bits_data_0_12(tensorStore_io_tensor_wr_bits_data_0_12),
    .io_tensor_wr_bits_data_0_13(tensorStore_io_tensor_wr_bits_data_0_13),
    .io_tensor_wr_bits_data_0_14(tensorStore_io_tensor_wr_bits_data_0_14),
    .io_tensor_wr_bits_data_0_15(tensorStore_io_tensor_wr_bits_data_0_15)
  );
  assign _T_597 = dec_io_pop_prev ? s_io_sready : 1'h1; // @[Store.scala 54:40:@24617.4]
  assign start = inst_q_io_deq_valid & _T_597; // @[Store.scala 54:35:@24618.4]
  assign _T_598 = 2'h0 == state; // @[Conditional.scala 37:30:@24619.4]
  assign _GEN_0 = dec_io_isStore ? 2'h2 : state; // @[Store.scala 63:36:@24626.10]
  assign _GEN_1 = dec_io_isSync ? 2'h1 : _GEN_0; // @[Store.scala 61:29:@24622.8]
  assign _GEN_2 = start ? _GEN_1 : state; // @[Store.scala 60:19:@24621.6]
  assign _T_599 = 2'h1 == state; // @[Conditional.scala 37:30:@24632.6]
  assign _T_600 = 2'h2 == state; // @[Conditional.scala 37:30:@24637.8]
  assign _GEN_3 = tensorStore_io_done ? 2'h0 : state; // @[Store.scala 72:18:@24639.10]
  assign _GEN_4 = _T_600 ? _GEN_3 : state; // @[Conditional.scala 39:67:@24638.8]
  assign _GEN_5 = _T_599 ? 2'h0 : _GEN_4; // @[Conditional.scala 39:67:@24633.6]
  assign _GEN_6 = _T_598 ? _GEN_2 : _GEN_5; // @[Conditional.scala 40:58:@24620.4]
  assign _T_601 = state == 2'h2; // @[Store.scala 80:33:@24646.4]
  assign _T_602 = _T_601 & tensorStore_io_done; // @[Store.scala 80:42:@24647.4]
  assign _T_603 = state == 2'h1; // @[Store.scala 80:59:@24648.4]
  assign _T_604 = _T_602 | _T_603; // @[Store.scala 80:50:@24649.4]
  assign _T_605 = state == 2'h0; // @[Store.scala 83:33:@24651.4]
  assign _T_606 = _T_605 & start; // @[Store.scala 83:43:@24652.4]
  assign io_o_post = dec_io_push_prev & _T_604; // @[Store.scala 92:13:@24712.4]
  assign io_inst_ready = inst_q_io_enq_ready; // @[Store.scala 79:17:@24645.4]
  assign io_vme_wr_cmd_valid = tensorStore_io_vme_wr_cmd_valid; // @[Store.scala 86:13:@24663.4]
  assign io_vme_wr_cmd_bits_addr = tensorStore_io_vme_wr_cmd_bits_addr; // @[Store.scala 86:13:@24662.4]
  assign io_vme_wr_cmd_bits_len = tensorStore_io_vme_wr_cmd_bits_len; // @[Store.scala 86:13:@24661.4]
  assign io_vme_wr_data_valid = tensorStore_io_vme_wr_data_valid; // @[Store.scala 86:13:@24659.4]
  assign io_vme_wr_data_bits = tensorStore_io_vme_wr_data_bits; // @[Store.scala 86:13:@24658.4]
  assign s_clock = clock; // @[:@24605.4]
  assign s_reset = reset; // @[:@24606.4]
  assign s_io_spost = io_i_post; // @[Store.scala 90:14:@24702.4]
  assign s_io_swait = dec_io_pop_prev & _T_606; // @[Store.scala 91:14:@24706.4]
  assign inst_q_clock = clock; // @[:@24608.4]
  assign inst_q_reset = reset; // @[:@24609.4]
  assign inst_q_io_enq_valid = io_inst_valid; // @[Store.scala 79:17:@24644.4]
  assign inst_q_io_enq_bits = io_inst_bits; // @[Store.scala 79:17:@24643.4]
  assign inst_q_io_deq_ready = _T_602 | _T_603; // @[Store.scala 80:23:@24650.4]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Store.scala 50:15:@24613.4]
  assign tensorStore_clock = clock; // @[:@24615.4]
  assign tensorStore_reset = reset; // @[:@24616.4]
  assign tensorStore_io_start = _T_606 & dec_io_isStore; // @[Store.scala 83:24:@24654.4]
  assign tensorStore_io_inst = inst_q_io_deq_bits; // @[Store.scala 84:23:@24655.4]
  assign tensorStore_io_baddr = io_out_baddr; // @[Store.scala 85:24:@24656.4]
  assign tensorStore_io_vme_wr_cmd_ready = io_vme_wr_cmd_ready; // @[Store.scala 86:13:@24664.4]
  assign tensorStore_io_vme_wr_data_ready = io_vme_wr_data_ready; // @[Store.scala 86:13:@24660.4]
  assign tensorStore_io_vme_wr_ack = io_vme_wr_ack; // @[Store.scala 86:13:@24657.4]
  assign tensorStore_io_tensor_wr_valid = io_out_wr_valid; // @[Store.scala 87:25:@24682.4]
  assign tensorStore_io_tensor_wr_bits_idx = io_out_wr_bits_idx; // @[Store.scala 87:25:@24681.4]
  assign tensorStore_io_tensor_wr_bits_data_0_0 = io_out_wr_bits_data_0_0; // @[Store.scala 87:25:@24665.4]
  assign tensorStore_io_tensor_wr_bits_data_0_1 = io_out_wr_bits_data_0_1; // @[Store.scala 87:25:@24666.4]
  assign tensorStore_io_tensor_wr_bits_data_0_2 = io_out_wr_bits_data_0_2; // @[Store.scala 87:25:@24667.4]
  assign tensorStore_io_tensor_wr_bits_data_0_3 = io_out_wr_bits_data_0_3; // @[Store.scala 87:25:@24668.4]
  assign tensorStore_io_tensor_wr_bits_data_0_4 = io_out_wr_bits_data_0_4; // @[Store.scala 87:25:@24669.4]
  assign tensorStore_io_tensor_wr_bits_data_0_5 = io_out_wr_bits_data_0_5; // @[Store.scala 87:25:@24670.4]
  assign tensorStore_io_tensor_wr_bits_data_0_6 = io_out_wr_bits_data_0_6; // @[Store.scala 87:25:@24671.4]
  assign tensorStore_io_tensor_wr_bits_data_0_7 = io_out_wr_bits_data_0_7; // @[Store.scala 87:25:@24672.4]
  assign tensorStore_io_tensor_wr_bits_data_0_8 = io_out_wr_bits_data_0_8; // @[Store.scala 87:25:@24673.4]
  assign tensorStore_io_tensor_wr_bits_data_0_9 = io_out_wr_bits_data_0_9; // @[Store.scala 87:25:@24674.4]
  assign tensorStore_io_tensor_wr_bits_data_0_10 = io_out_wr_bits_data_0_10; // @[Store.scala 87:25:@24675.4]
  assign tensorStore_io_tensor_wr_bits_data_0_11 = io_out_wr_bits_data_0_11; // @[Store.scala 87:25:@24676.4]
  assign tensorStore_io_tensor_wr_bits_data_0_12 = io_out_wr_bits_data_0_12; // @[Store.scala 87:25:@24677.4]
  assign tensorStore_io_tensor_wr_bits_data_0_13 = io_out_wr_bits_data_0_13; // @[Store.scala 87:25:@24678.4]
  assign tensorStore_io_tensor_wr_bits_data_0_14 = io_out_wr_bits_data_0_14; // @[Store.scala 87:25:@24679.4]
  assign tensorStore_io_tensor_wr_bits_data_0_15 = io_out_wr_bits_data_0_15; // @[Store.scala 87:25:@24680.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_598) begin
        if (start) begin
          if (dec_io_isSync) begin
            state <= 2'h1;
          end else begin
            if (dec_io_isStore) begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_599) begin
          state <= 2'h0;
        end else begin
          if (_T_600) begin
            if (tensorStore_io_done) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module EventCounters( // @[:@24714.2]
  input         clock, // @[:@24715.4]
  input         reset, // @[:@24716.4]
  input         io_launch, // @[:@24717.4]
  input         io_finish, // @[:@24717.4]
  output        io_ecnt_0_valid, // @[:@24717.4]
  output [31:0] io_ecnt_0_bits, // @[:@24717.4]
  output        io_ucnt_0_valid, // @[:@24717.4]
  output [31:0] io_ucnt_0_bits, // @[:@24717.4]
  input         io_acc_wr_event // @[:@24717.4]
);
  reg [31:0] cycle_cnt; // @[EventCounters.scala 50:26:@24719.4]
  reg [31:0] _RAND_0;
  wire  _T_38; // @[EventCounters.scala 51:21:@24720.4]
  wire  _T_39; // @[EventCounters.scala 51:18:@24721.4]
  wire [32:0] _T_41; // @[EventCounters.scala 52:28:@24723.6]
  wire [31:0] _T_42; // @[EventCounters.scala 52:28:@24724.6]
  wire [31:0] _GEN_0; // @[EventCounters.scala 51:33:@24722.4]
  reg [31:0] acc_wr_count; // @[EventCounters.scala 59:25:@24732.4]
  reg [31:0] _RAND_1;
  wire  _T_46; // @[EventCounters.scala 60:9:@24733.4]
  wire  _T_47; // @[EventCounters.scala 60:20:@24734.4]
  wire [32:0] _T_50; // @[EventCounters.scala 63:34:@24740.8]
  wire [31:0] _T_51; // @[EventCounters.scala 63:34:@24741.8]
  wire [31:0] _GEN_1; // @[EventCounters.scala 62:32:@24739.6]
  assign _T_38 = io_finish == 1'h0; // @[EventCounters.scala 51:21:@24720.4]
  assign _T_39 = io_launch & _T_38; // @[EventCounters.scala 51:18:@24721.4]
  assign _T_41 = cycle_cnt + 32'h1; // @[EventCounters.scala 52:28:@24723.6]
  assign _T_42 = cycle_cnt + 32'h1; // @[EventCounters.scala 52:28:@24724.6]
  assign _GEN_0 = _T_39 ? _T_42 : 32'h0; // @[EventCounters.scala 51:33:@24722.4]
  assign _T_46 = io_launch == 1'h0; // @[EventCounters.scala 60:9:@24733.4]
  assign _T_47 = _T_46 | io_finish; // @[EventCounters.scala 60:20:@24734.4]
  assign _T_50 = acc_wr_count + 32'h1; // @[EventCounters.scala 63:34:@24740.8]
  assign _T_51 = acc_wr_count + 32'h1; // @[EventCounters.scala 63:34:@24741.8]
  assign _GEN_1 = io_acc_wr_event ? _T_51 : acc_wr_count; // @[EventCounters.scala 62:32:@24739.6]
  assign io_ecnt_0_valid = io_finish; // @[EventCounters.scala 56:20:@24730.4]
  assign io_ecnt_0_bits = cycle_cnt; // @[EventCounters.scala 57:19:@24731.4]
  assign io_ucnt_0_valid = io_finish; // @[EventCounters.scala 65:20:@24744.4]
  assign io_ucnt_0_bits = acc_wr_count; // @[EventCounters.scala 66:19:@24745.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycle_cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  acc_wr_count = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cycle_cnt <= 32'h0;
    end else begin
      if (_T_39) begin
        cycle_cnt <= _T_42;
      end else begin
        cycle_cnt <= 32'h0;
      end
    end
    if (_T_47) begin
      acc_wr_count <= 32'h0;
    end else begin
      if (io_acc_wr_event) begin
        acc_wr_count <= _T_51;
      end
    end
  end
endmodule
module Core( // @[:@24747.2]
  input         clock, // @[:@24748.4]
  input         reset, // @[:@24749.4]
  input         io_vcr_launch, // @[:@24750.4]
  output        io_vcr_finish, // @[:@24750.4]
  output        io_vcr_ecnt_0_valid, // @[:@24750.4]
  output [31:0] io_vcr_ecnt_0_bits, // @[:@24750.4]
  input  [31:0] io_vcr_vals_0, // @[:@24750.4]
  input  [31:0] io_vcr_ptrs_0, // @[:@24750.4]
  input  [31:0] io_vcr_ptrs_1, // @[:@24750.4]
  input  [31:0] io_vcr_ptrs_2, // @[:@24750.4]
  input  [31:0] io_vcr_ptrs_3, // @[:@24750.4]
  input  [31:0] io_vcr_ptrs_4, // @[:@24750.4]
  input  [31:0] io_vcr_ptrs_5, // @[:@24750.4]
  output        io_vcr_ucnt_0_valid, // @[:@24750.4]
  output [31:0] io_vcr_ucnt_0_bits, // @[:@24750.4]
  input         io_vme_rd_0_cmd_ready, // @[:@24750.4]
  output        io_vme_rd_0_cmd_valid, // @[:@24750.4]
  output [31:0] io_vme_rd_0_cmd_bits_addr, // @[:@24750.4]
  output [7:0]  io_vme_rd_0_cmd_bits_len, // @[:@24750.4]
  output        io_vme_rd_0_data_ready, // @[:@24750.4]
  input         io_vme_rd_0_data_valid, // @[:@24750.4]
  input  [63:0] io_vme_rd_0_data_bits, // @[:@24750.4]
  input         io_vme_rd_1_cmd_ready, // @[:@24750.4]
  output        io_vme_rd_1_cmd_valid, // @[:@24750.4]
  output [31:0] io_vme_rd_1_cmd_bits_addr, // @[:@24750.4]
  output [7:0]  io_vme_rd_1_cmd_bits_len, // @[:@24750.4]
  output        io_vme_rd_1_data_ready, // @[:@24750.4]
  input         io_vme_rd_1_data_valid, // @[:@24750.4]
  input  [63:0] io_vme_rd_1_data_bits, // @[:@24750.4]
  input         io_vme_rd_2_cmd_ready, // @[:@24750.4]
  output        io_vme_rd_2_cmd_valid, // @[:@24750.4]
  output [31:0] io_vme_rd_2_cmd_bits_addr, // @[:@24750.4]
  output [7:0]  io_vme_rd_2_cmd_bits_len, // @[:@24750.4]
  output        io_vme_rd_2_data_ready, // @[:@24750.4]
  input         io_vme_rd_2_data_valid, // @[:@24750.4]
  input  [63:0] io_vme_rd_2_data_bits, // @[:@24750.4]
  input         io_vme_rd_3_cmd_ready, // @[:@24750.4]
  output        io_vme_rd_3_cmd_valid, // @[:@24750.4]
  output [31:0] io_vme_rd_3_cmd_bits_addr, // @[:@24750.4]
  output [7:0]  io_vme_rd_3_cmd_bits_len, // @[:@24750.4]
  output        io_vme_rd_3_data_ready, // @[:@24750.4]
  input         io_vme_rd_3_data_valid, // @[:@24750.4]
  input  [63:0] io_vme_rd_3_data_bits, // @[:@24750.4]
  input         io_vme_rd_4_cmd_ready, // @[:@24750.4]
  output        io_vme_rd_4_cmd_valid, // @[:@24750.4]
  output [31:0] io_vme_rd_4_cmd_bits_addr, // @[:@24750.4]
  output [7:0]  io_vme_rd_4_cmd_bits_len, // @[:@24750.4]
  output        io_vme_rd_4_data_ready, // @[:@24750.4]
  input         io_vme_rd_4_data_valid, // @[:@24750.4]
  input  [63:0] io_vme_rd_4_data_bits, // @[:@24750.4]
  input         io_vme_wr_0_cmd_ready, // @[:@24750.4]
  output        io_vme_wr_0_cmd_valid, // @[:@24750.4]
  output [31:0] io_vme_wr_0_cmd_bits_addr, // @[:@24750.4]
  output [7:0]  io_vme_wr_0_cmd_bits_len, // @[:@24750.4]
  input         io_vme_wr_0_data_ready, // @[:@24750.4]
  output        io_vme_wr_0_data_valid, // @[:@24750.4]
  output [63:0] io_vme_wr_0_data_bits, // @[:@24750.4]
  input         io_vme_wr_0_ack // @[:@24750.4]
);
  wire  fetch_clock; // @[Core.scala 66:21:@24752.4]
  wire  fetch_reset; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_launch; // @[Core.scala 66:21:@24752.4]
  wire [31:0] fetch_io_ins_baddr; // @[Core.scala 66:21:@24752.4]
  wire [31:0] fetch_io_ins_count; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_vme_rd_cmd_ready; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_vme_rd_cmd_valid; // @[Core.scala 66:21:@24752.4]
  wire [31:0] fetch_io_vme_rd_cmd_bits_addr; // @[Core.scala 66:21:@24752.4]
  wire [7:0] fetch_io_vme_rd_cmd_bits_len; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_vme_rd_data_ready; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_vme_rd_data_valid; // @[Core.scala 66:21:@24752.4]
  wire [63:0] fetch_io_vme_rd_data_bits; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_inst_ld_ready; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_inst_ld_valid; // @[Core.scala 66:21:@24752.4]
  wire [127:0] fetch_io_inst_ld_bits; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_inst_co_ready; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_inst_co_valid; // @[Core.scala 66:21:@24752.4]
  wire [127:0] fetch_io_inst_co_bits; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_inst_st_ready; // @[Core.scala 66:21:@24752.4]
  wire  fetch_io_inst_st_valid; // @[Core.scala 66:21:@24752.4]
  wire [127:0] fetch_io_inst_st_bits; // @[Core.scala 66:21:@24752.4]
  wire  load_clock; // @[Core.scala 67:20:@24755.4]
  wire  load_reset; // @[Core.scala 67:20:@24755.4]
  wire  load_io_i_post; // @[Core.scala 67:20:@24755.4]
  wire  load_io_o_post; // @[Core.scala 67:20:@24755.4]
  wire  load_io_inst_ready; // @[Core.scala 67:20:@24755.4]
  wire  load_io_inst_valid; // @[Core.scala 67:20:@24755.4]
  wire [127:0] load_io_inst_bits; // @[Core.scala 67:20:@24755.4]
  wire [31:0] load_io_inp_baddr; // @[Core.scala 67:20:@24755.4]
  wire [31:0] load_io_wgt_baddr; // @[Core.scala 67:20:@24755.4]
  wire  load_io_vme_rd_0_cmd_ready; // @[Core.scala 67:20:@24755.4]
  wire  load_io_vme_rd_0_cmd_valid; // @[Core.scala 67:20:@24755.4]
  wire [31:0] load_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_vme_rd_0_cmd_bits_len; // @[Core.scala 67:20:@24755.4]
  wire  load_io_vme_rd_0_data_ready; // @[Core.scala 67:20:@24755.4]
  wire  load_io_vme_rd_0_data_valid; // @[Core.scala 67:20:@24755.4]
  wire [63:0] load_io_vme_rd_0_data_bits; // @[Core.scala 67:20:@24755.4]
  wire  load_io_vme_rd_1_cmd_ready; // @[Core.scala 67:20:@24755.4]
  wire  load_io_vme_rd_1_cmd_valid; // @[Core.scala 67:20:@24755.4]
  wire [31:0] load_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_vme_rd_1_cmd_bits_len; // @[Core.scala 67:20:@24755.4]
  wire  load_io_vme_rd_1_data_ready; // @[Core.scala 67:20:@24755.4]
  wire  load_io_vme_rd_1_data_valid; // @[Core.scala 67:20:@24755.4]
  wire [63:0] load_io_vme_rd_1_data_bits; // @[Core.scala 67:20:@24755.4]
  wire  load_io_inp_rd_idx_valid; // @[Core.scala 67:20:@24755.4]
  wire [10:0] load_io_inp_rd_idx_bits; // @[Core.scala 67:20:@24755.4]
  wire  load_io_inp_rd_data_valid; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_inp_rd_data_bits_0_15; // @[Core.scala 67:20:@24755.4]
  wire  load_io_wgt_rd_idx_valid; // @[Core.scala 67:20:@24755.4]
  wire [9:0] load_io_wgt_rd_idx_bits; // @[Core.scala 67:20:@24755.4]
  wire  load_io_wgt_rd_data_valid; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_0_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_1_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_2_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_3_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_4_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_5_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_6_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_7_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_8_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_9_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_10_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_11_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_12_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_13_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_14_15; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_0; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_1; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_2; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_3; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_4; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_5; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_6; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_7; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_8; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_9; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_10; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_11; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_12; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_13; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_14; // @[Core.scala 67:20:@24755.4]
  wire [7:0] load_io_wgt_rd_data_bits_15_15; // @[Core.scala 67:20:@24755.4]
  wire  compute_clock; // @[Core.scala 68:23:@24758.4]
  wire  compute_reset; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_i_post_0; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_i_post_1; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_o_post_0; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_o_post_1; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_inst_ready; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_inst_valid; // @[Core.scala 68:23:@24758.4]
  wire [127:0] compute_io_inst_bits; // @[Core.scala 68:23:@24758.4]
  wire [31:0] compute_io_uop_baddr; // @[Core.scala 68:23:@24758.4]
  wire [31:0] compute_io_acc_baddr; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_vme_rd_0_cmd_ready; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_vme_rd_0_cmd_valid; // @[Core.scala 68:23:@24758.4]
  wire [31:0] compute_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_vme_rd_0_cmd_bits_len; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_vme_rd_0_data_ready; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_vme_rd_0_data_valid; // @[Core.scala 68:23:@24758.4]
  wire [63:0] compute_io_vme_rd_0_data_bits; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_vme_rd_1_cmd_ready; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_vme_rd_1_cmd_valid; // @[Core.scala 68:23:@24758.4]
  wire [31:0] compute_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_vme_rd_1_cmd_bits_len; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_vme_rd_1_data_ready; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_vme_rd_1_data_valid; // @[Core.scala 68:23:@24758.4]
  wire [63:0] compute_io_vme_rd_1_data_bits; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_inp_rd_idx_valid; // @[Core.scala 68:23:@24758.4]
  wire [10:0] compute_io_inp_rd_idx_bits; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_inp_rd_data_valid; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_inp_rd_data_bits_0_15; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_wgt_rd_idx_valid; // @[Core.scala 68:23:@24758.4]
  wire [9:0] compute_io_wgt_rd_idx_bits; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_wgt_rd_data_valid; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_0_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_1_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_2_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_3_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_4_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_5_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_6_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_7_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_8_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_9_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_10_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_11_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_12_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_13_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_14_15; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_wgt_rd_data_bits_15_15; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_out_wr_valid; // @[Core.scala 68:23:@24758.4]
  wire [10:0] compute_io_out_wr_bits_idx; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_0; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_1; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_2; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_3; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_4; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_5; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_6; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_7; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_8; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_9; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_10; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_11; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_12; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_13; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_14; // @[Core.scala 68:23:@24758.4]
  wire [7:0] compute_io_out_wr_bits_data_0_15; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_finish; // @[Core.scala 68:23:@24758.4]
  wire  compute_io_acc_wr_event; // @[Core.scala 68:23:@24758.4]
  wire  store_clock; // @[Core.scala 69:21:@24761.4]
  wire  store_reset; // @[Core.scala 69:21:@24761.4]
  wire  store_io_i_post; // @[Core.scala 69:21:@24761.4]
  wire  store_io_o_post; // @[Core.scala 69:21:@24761.4]
  wire  store_io_inst_ready; // @[Core.scala 69:21:@24761.4]
  wire  store_io_inst_valid; // @[Core.scala 69:21:@24761.4]
  wire [127:0] store_io_inst_bits; // @[Core.scala 69:21:@24761.4]
  wire [31:0] store_io_out_baddr; // @[Core.scala 69:21:@24761.4]
  wire  store_io_vme_wr_cmd_ready; // @[Core.scala 69:21:@24761.4]
  wire  store_io_vme_wr_cmd_valid; // @[Core.scala 69:21:@24761.4]
  wire [31:0] store_io_vme_wr_cmd_bits_addr; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_vme_wr_cmd_bits_len; // @[Core.scala 69:21:@24761.4]
  wire  store_io_vme_wr_data_ready; // @[Core.scala 69:21:@24761.4]
  wire  store_io_vme_wr_data_valid; // @[Core.scala 69:21:@24761.4]
  wire [63:0] store_io_vme_wr_data_bits; // @[Core.scala 69:21:@24761.4]
  wire  store_io_vme_wr_ack; // @[Core.scala 69:21:@24761.4]
  wire  store_io_out_wr_valid; // @[Core.scala 69:21:@24761.4]
  wire [10:0] store_io_out_wr_bits_idx; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_0; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_1; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_2; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_3; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_4; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_5; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_6; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_7; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_8; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_9; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_10; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_11; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_12; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_13; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_14; // @[Core.scala 69:21:@24761.4]
  wire [7:0] store_io_out_wr_bits_data_0_15; // @[Core.scala 69:21:@24761.4]
  wire  ecounters_clock; // @[Core.scala 70:25:@24764.4]
  wire  ecounters_reset; // @[Core.scala 70:25:@24764.4]
  wire  ecounters_io_launch; // @[Core.scala 70:25:@24764.4]
  wire  ecounters_io_finish; // @[Core.scala 70:25:@24764.4]
  wire  ecounters_io_ecnt_0_valid; // @[Core.scala 70:25:@24764.4]
  wire [31:0] ecounters_io_ecnt_0_bits; // @[Core.scala 70:25:@24764.4]
  wire  ecounters_io_ucnt_0_valid; // @[Core.scala 70:25:@24764.4]
  wire [31:0] ecounters_io_ucnt_0_bits; // @[Core.scala 70:25:@24764.4]
  wire  ecounters_io_acc_wr_event; // @[Core.scala 70:25:@24764.4]
  reg  finish; // @[Core.scala 118:23:@25429.4]
  reg [31:0] _RAND_0;
  Fetch fetch ( // @[Core.scala 66:21:@24752.4]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_launch(fetch_io_launch),
    .io_ins_baddr(fetch_io_ins_baddr),
    .io_ins_count(fetch_io_ins_count),
    .io_vme_rd_cmd_ready(fetch_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(fetch_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(fetch_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(fetch_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(fetch_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(fetch_io_vme_rd_data_valid),
    .io_vme_rd_data_bits(fetch_io_vme_rd_data_bits),
    .io_inst_ld_ready(fetch_io_inst_ld_ready),
    .io_inst_ld_valid(fetch_io_inst_ld_valid),
    .io_inst_ld_bits(fetch_io_inst_ld_bits),
    .io_inst_co_ready(fetch_io_inst_co_ready),
    .io_inst_co_valid(fetch_io_inst_co_valid),
    .io_inst_co_bits(fetch_io_inst_co_bits),
    .io_inst_st_ready(fetch_io_inst_st_ready),
    .io_inst_st_valid(fetch_io_inst_st_valid),
    .io_inst_st_bits(fetch_io_inst_st_bits)
  );
  Load load ( // @[Core.scala 67:20:@24755.4]
    .clock(load_clock),
    .reset(load_reset),
    .io_i_post(load_io_i_post),
    .io_o_post(load_io_o_post),
    .io_inst_ready(load_io_inst_ready),
    .io_inst_valid(load_io_inst_valid),
    .io_inst_bits(load_io_inst_bits),
    .io_inp_baddr(load_io_inp_baddr),
    .io_wgt_baddr(load_io_wgt_baddr),
    .io_vme_rd_0_cmd_ready(load_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(load_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(load_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(load_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(load_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(load_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits(load_io_vme_rd_0_data_bits),
    .io_vme_rd_1_cmd_ready(load_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(load_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(load_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(load_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_data_ready(load_io_vme_rd_1_data_ready),
    .io_vme_rd_1_data_valid(load_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits(load_io_vme_rd_1_data_bits),
    .io_inp_rd_idx_valid(load_io_inp_rd_idx_valid),
    .io_inp_rd_idx_bits(load_io_inp_rd_idx_bits),
    .io_inp_rd_data_valid(load_io_inp_rd_data_valid),
    .io_inp_rd_data_bits_0_0(load_io_inp_rd_data_bits_0_0),
    .io_inp_rd_data_bits_0_1(load_io_inp_rd_data_bits_0_1),
    .io_inp_rd_data_bits_0_2(load_io_inp_rd_data_bits_0_2),
    .io_inp_rd_data_bits_0_3(load_io_inp_rd_data_bits_0_3),
    .io_inp_rd_data_bits_0_4(load_io_inp_rd_data_bits_0_4),
    .io_inp_rd_data_bits_0_5(load_io_inp_rd_data_bits_0_5),
    .io_inp_rd_data_bits_0_6(load_io_inp_rd_data_bits_0_6),
    .io_inp_rd_data_bits_0_7(load_io_inp_rd_data_bits_0_7),
    .io_inp_rd_data_bits_0_8(load_io_inp_rd_data_bits_0_8),
    .io_inp_rd_data_bits_0_9(load_io_inp_rd_data_bits_0_9),
    .io_inp_rd_data_bits_0_10(load_io_inp_rd_data_bits_0_10),
    .io_inp_rd_data_bits_0_11(load_io_inp_rd_data_bits_0_11),
    .io_inp_rd_data_bits_0_12(load_io_inp_rd_data_bits_0_12),
    .io_inp_rd_data_bits_0_13(load_io_inp_rd_data_bits_0_13),
    .io_inp_rd_data_bits_0_14(load_io_inp_rd_data_bits_0_14),
    .io_inp_rd_data_bits_0_15(load_io_inp_rd_data_bits_0_15),
    .io_wgt_rd_idx_valid(load_io_wgt_rd_idx_valid),
    .io_wgt_rd_idx_bits(load_io_wgt_rd_idx_bits),
    .io_wgt_rd_data_valid(load_io_wgt_rd_data_valid),
    .io_wgt_rd_data_bits_0_0(load_io_wgt_rd_data_bits_0_0),
    .io_wgt_rd_data_bits_0_1(load_io_wgt_rd_data_bits_0_1),
    .io_wgt_rd_data_bits_0_2(load_io_wgt_rd_data_bits_0_2),
    .io_wgt_rd_data_bits_0_3(load_io_wgt_rd_data_bits_0_3),
    .io_wgt_rd_data_bits_0_4(load_io_wgt_rd_data_bits_0_4),
    .io_wgt_rd_data_bits_0_5(load_io_wgt_rd_data_bits_0_5),
    .io_wgt_rd_data_bits_0_6(load_io_wgt_rd_data_bits_0_6),
    .io_wgt_rd_data_bits_0_7(load_io_wgt_rd_data_bits_0_7),
    .io_wgt_rd_data_bits_0_8(load_io_wgt_rd_data_bits_0_8),
    .io_wgt_rd_data_bits_0_9(load_io_wgt_rd_data_bits_0_9),
    .io_wgt_rd_data_bits_0_10(load_io_wgt_rd_data_bits_0_10),
    .io_wgt_rd_data_bits_0_11(load_io_wgt_rd_data_bits_0_11),
    .io_wgt_rd_data_bits_0_12(load_io_wgt_rd_data_bits_0_12),
    .io_wgt_rd_data_bits_0_13(load_io_wgt_rd_data_bits_0_13),
    .io_wgt_rd_data_bits_0_14(load_io_wgt_rd_data_bits_0_14),
    .io_wgt_rd_data_bits_0_15(load_io_wgt_rd_data_bits_0_15),
    .io_wgt_rd_data_bits_1_0(load_io_wgt_rd_data_bits_1_0),
    .io_wgt_rd_data_bits_1_1(load_io_wgt_rd_data_bits_1_1),
    .io_wgt_rd_data_bits_1_2(load_io_wgt_rd_data_bits_1_2),
    .io_wgt_rd_data_bits_1_3(load_io_wgt_rd_data_bits_1_3),
    .io_wgt_rd_data_bits_1_4(load_io_wgt_rd_data_bits_1_4),
    .io_wgt_rd_data_bits_1_5(load_io_wgt_rd_data_bits_1_5),
    .io_wgt_rd_data_bits_1_6(load_io_wgt_rd_data_bits_1_6),
    .io_wgt_rd_data_bits_1_7(load_io_wgt_rd_data_bits_1_7),
    .io_wgt_rd_data_bits_1_8(load_io_wgt_rd_data_bits_1_8),
    .io_wgt_rd_data_bits_1_9(load_io_wgt_rd_data_bits_1_9),
    .io_wgt_rd_data_bits_1_10(load_io_wgt_rd_data_bits_1_10),
    .io_wgt_rd_data_bits_1_11(load_io_wgt_rd_data_bits_1_11),
    .io_wgt_rd_data_bits_1_12(load_io_wgt_rd_data_bits_1_12),
    .io_wgt_rd_data_bits_1_13(load_io_wgt_rd_data_bits_1_13),
    .io_wgt_rd_data_bits_1_14(load_io_wgt_rd_data_bits_1_14),
    .io_wgt_rd_data_bits_1_15(load_io_wgt_rd_data_bits_1_15),
    .io_wgt_rd_data_bits_2_0(load_io_wgt_rd_data_bits_2_0),
    .io_wgt_rd_data_bits_2_1(load_io_wgt_rd_data_bits_2_1),
    .io_wgt_rd_data_bits_2_2(load_io_wgt_rd_data_bits_2_2),
    .io_wgt_rd_data_bits_2_3(load_io_wgt_rd_data_bits_2_3),
    .io_wgt_rd_data_bits_2_4(load_io_wgt_rd_data_bits_2_4),
    .io_wgt_rd_data_bits_2_5(load_io_wgt_rd_data_bits_2_5),
    .io_wgt_rd_data_bits_2_6(load_io_wgt_rd_data_bits_2_6),
    .io_wgt_rd_data_bits_2_7(load_io_wgt_rd_data_bits_2_7),
    .io_wgt_rd_data_bits_2_8(load_io_wgt_rd_data_bits_2_8),
    .io_wgt_rd_data_bits_2_9(load_io_wgt_rd_data_bits_2_9),
    .io_wgt_rd_data_bits_2_10(load_io_wgt_rd_data_bits_2_10),
    .io_wgt_rd_data_bits_2_11(load_io_wgt_rd_data_bits_2_11),
    .io_wgt_rd_data_bits_2_12(load_io_wgt_rd_data_bits_2_12),
    .io_wgt_rd_data_bits_2_13(load_io_wgt_rd_data_bits_2_13),
    .io_wgt_rd_data_bits_2_14(load_io_wgt_rd_data_bits_2_14),
    .io_wgt_rd_data_bits_2_15(load_io_wgt_rd_data_bits_2_15),
    .io_wgt_rd_data_bits_3_0(load_io_wgt_rd_data_bits_3_0),
    .io_wgt_rd_data_bits_3_1(load_io_wgt_rd_data_bits_3_1),
    .io_wgt_rd_data_bits_3_2(load_io_wgt_rd_data_bits_3_2),
    .io_wgt_rd_data_bits_3_3(load_io_wgt_rd_data_bits_3_3),
    .io_wgt_rd_data_bits_3_4(load_io_wgt_rd_data_bits_3_4),
    .io_wgt_rd_data_bits_3_5(load_io_wgt_rd_data_bits_3_5),
    .io_wgt_rd_data_bits_3_6(load_io_wgt_rd_data_bits_3_6),
    .io_wgt_rd_data_bits_3_7(load_io_wgt_rd_data_bits_3_7),
    .io_wgt_rd_data_bits_3_8(load_io_wgt_rd_data_bits_3_8),
    .io_wgt_rd_data_bits_3_9(load_io_wgt_rd_data_bits_3_9),
    .io_wgt_rd_data_bits_3_10(load_io_wgt_rd_data_bits_3_10),
    .io_wgt_rd_data_bits_3_11(load_io_wgt_rd_data_bits_3_11),
    .io_wgt_rd_data_bits_3_12(load_io_wgt_rd_data_bits_3_12),
    .io_wgt_rd_data_bits_3_13(load_io_wgt_rd_data_bits_3_13),
    .io_wgt_rd_data_bits_3_14(load_io_wgt_rd_data_bits_3_14),
    .io_wgt_rd_data_bits_3_15(load_io_wgt_rd_data_bits_3_15),
    .io_wgt_rd_data_bits_4_0(load_io_wgt_rd_data_bits_4_0),
    .io_wgt_rd_data_bits_4_1(load_io_wgt_rd_data_bits_4_1),
    .io_wgt_rd_data_bits_4_2(load_io_wgt_rd_data_bits_4_2),
    .io_wgt_rd_data_bits_4_3(load_io_wgt_rd_data_bits_4_3),
    .io_wgt_rd_data_bits_4_4(load_io_wgt_rd_data_bits_4_4),
    .io_wgt_rd_data_bits_4_5(load_io_wgt_rd_data_bits_4_5),
    .io_wgt_rd_data_bits_4_6(load_io_wgt_rd_data_bits_4_6),
    .io_wgt_rd_data_bits_4_7(load_io_wgt_rd_data_bits_4_7),
    .io_wgt_rd_data_bits_4_8(load_io_wgt_rd_data_bits_4_8),
    .io_wgt_rd_data_bits_4_9(load_io_wgt_rd_data_bits_4_9),
    .io_wgt_rd_data_bits_4_10(load_io_wgt_rd_data_bits_4_10),
    .io_wgt_rd_data_bits_4_11(load_io_wgt_rd_data_bits_4_11),
    .io_wgt_rd_data_bits_4_12(load_io_wgt_rd_data_bits_4_12),
    .io_wgt_rd_data_bits_4_13(load_io_wgt_rd_data_bits_4_13),
    .io_wgt_rd_data_bits_4_14(load_io_wgt_rd_data_bits_4_14),
    .io_wgt_rd_data_bits_4_15(load_io_wgt_rd_data_bits_4_15),
    .io_wgt_rd_data_bits_5_0(load_io_wgt_rd_data_bits_5_0),
    .io_wgt_rd_data_bits_5_1(load_io_wgt_rd_data_bits_5_1),
    .io_wgt_rd_data_bits_5_2(load_io_wgt_rd_data_bits_5_2),
    .io_wgt_rd_data_bits_5_3(load_io_wgt_rd_data_bits_5_3),
    .io_wgt_rd_data_bits_5_4(load_io_wgt_rd_data_bits_5_4),
    .io_wgt_rd_data_bits_5_5(load_io_wgt_rd_data_bits_5_5),
    .io_wgt_rd_data_bits_5_6(load_io_wgt_rd_data_bits_5_6),
    .io_wgt_rd_data_bits_5_7(load_io_wgt_rd_data_bits_5_7),
    .io_wgt_rd_data_bits_5_8(load_io_wgt_rd_data_bits_5_8),
    .io_wgt_rd_data_bits_5_9(load_io_wgt_rd_data_bits_5_9),
    .io_wgt_rd_data_bits_5_10(load_io_wgt_rd_data_bits_5_10),
    .io_wgt_rd_data_bits_5_11(load_io_wgt_rd_data_bits_5_11),
    .io_wgt_rd_data_bits_5_12(load_io_wgt_rd_data_bits_5_12),
    .io_wgt_rd_data_bits_5_13(load_io_wgt_rd_data_bits_5_13),
    .io_wgt_rd_data_bits_5_14(load_io_wgt_rd_data_bits_5_14),
    .io_wgt_rd_data_bits_5_15(load_io_wgt_rd_data_bits_5_15),
    .io_wgt_rd_data_bits_6_0(load_io_wgt_rd_data_bits_6_0),
    .io_wgt_rd_data_bits_6_1(load_io_wgt_rd_data_bits_6_1),
    .io_wgt_rd_data_bits_6_2(load_io_wgt_rd_data_bits_6_2),
    .io_wgt_rd_data_bits_6_3(load_io_wgt_rd_data_bits_6_3),
    .io_wgt_rd_data_bits_6_4(load_io_wgt_rd_data_bits_6_4),
    .io_wgt_rd_data_bits_6_5(load_io_wgt_rd_data_bits_6_5),
    .io_wgt_rd_data_bits_6_6(load_io_wgt_rd_data_bits_6_6),
    .io_wgt_rd_data_bits_6_7(load_io_wgt_rd_data_bits_6_7),
    .io_wgt_rd_data_bits_6_8(load_io_wgt_rd_data_bits_6_8),
    .io_wgt_rd_data_bits_6_9(load_io_wgt_rd_data_bits_6_9),
    .io_wgt_rd_data_bits_6_10(load_io_wgt_rd_data_bits_6_10),
    .io_wgt_rd_data_bits_6_11(load_io_wgt_rd_data_bits_6_11),
    .io_wgt_rd_data_bits_6_12(load_io_wgt_rd_data_bits_6_12),
    .io_wgt_rd_data_bits_6_13(load_io_wgt_rd_data_bits_6_13),
    .io_wgt_rd_data_bits_6_14(load_io_wgt_rd_data_bits_6_14),
    .io_wgt_rd_data_bits_6_15(load_io_wgt_rd_data_bits_6_15),
    .io_wgt_rd_data_bits_7_0(load_io_wgt_rd_data_bits_7_0),
    .io_wgt_rd_data_bits_7_1(load_io_wgt_rd_data_bits_7_1),
    .io_wgt_rd_data_bits_7_2(load_io_wgt_rd_data_bits_7_2),
    .io_wgt_rd_data_bits_7_3(load_io_wgt_rd_data_bits_7_3),
    .io_wgt_rd_data_bits_7_4(load_io_wgt_rd_data_bits_7_4),
    .io_wgt_rd_data_bits_7_5(load_io_wgt_rd_data_bits_7_5),
    .io_wgt_rd_data_bits_7_6(load_io_wgt_rd_data_bits_7_6),
    .io_wgt_rd_data_bits_7_7(load_io_wgt_rd_data_bits_7_7),
    .io_wgt_rd_data_bits_7_8(load_io_wgt_rd_data_bits_7_8),
    .io_wgt_rd_data_bits_7_9(load_io_wgt_rd_data_bits_7_9),
    .io_wgt_rd_data_bits_7_10(load_io_wgt_rd_data_bits_7_10),
    .io_wgt_rd_data_bits_7_11(load_io_wgt_rd_data_bits_7_11),
    .io_wgt_rd_data_bits_7_12(load_io_wgt_rd_data_bits_7_12),
    .io_wgt_rd_data_bits_7_13(load_io_wgt_rd_data_bits_7_13),
    .io_wgt_rd_data_bits_7_14(load_io_wgt_rd_data_bits_7_14),
    .io_wgt_rd_data_bits_7_15(load_io_wgt_rd_data_bits_7_15),
    .io_wgt_rd_data_bits_8_0(load_io_wgt_rd_data_bits_8_0),
    .io_wgt_rd_data_bits_8_1(load_io_wgt_rd_data_bits_8_1),
    .io_wgt_rd_data_bits_8_2(load_io_wgt_rd_data_bits_8_2),
    .io_wgt_rd_data_bits_8_3(load_io_wgt_rd_data_bits_8_3),
    .io_wgt_rd_data_bits_8_4(load_io_wgt_rd_data_bits_8_4),
    .io_wgt_rd_data_bits_8_5(load_io_wgt_rd_data_bits_8_5),
    .io_wgt_rd_data_bits_8_6(load_io_wgt_rd_data_bits_8_6),
    .io_wgt_rd_data_bits_8_7(load_io_wgt_rd_data_bits_8_7),
    .io_wgt_rd_data_bits_8_8(load_io_wgt_rd_data_bits_8_8),
    .io_wgt_rd_data_bits_8_9(load_io_wgt_rd_data_bits_8_9),
    .io_wgt_rd_data_bits_8_10(load_io_wgt_rd_data_bits_8_10),
    .io_wgt_rd_data_bits_8_11(load_io_wgt_rd_data_bits_8_11),
    .io_wgt_rd_data_bits_8_12(load_io_wgt_rd_data_bits_8_12),
    .io_wgt_rd_data_bits_8_13(load_io_wgt_rd_data_bits_8_13),
    .io_wgt_rd_data_bits_8_14(load_io_wgt_rd_data_bits_8_14),
    .io_wgt_rd_data_bits_8_15(load_io_wgt_rd_data_bits_8_15),
    .io_wgt_rd_data_bits_9_0(load_io_wgt_rd_data_bits_9_0),
    .io_wgt_rd_data_bits_9_1(load_io_wgt_rd_data_bits_9_1),
    .io_wgt_rd_data_bits_9_2(load_io_wgt_rd_data_bits_9_2),
    .io_wgt_rd_data_bits_9_3(load_io_wgt_rd_data_bits_9_3),
    .io_wgt_rd_data_bits_9_4(load_io_wgt_rd_data_bits_9_4),
    .io_wgt_rd_data_bits_9_5(load_io_wgt_rd_data_bits_9_5),
    .io_wgt_rd_data_bits_9_6(load_io_wgt_rd_data_bits_9_6),
    .io_wgt_rd_data_bits_9_7(load_io_wgt_rd_data_bits_9_7),
    .io_wgt_rd_data_bits_9_8(load_io_wgt_rd_data_bits_9_8),
    .io_wgt_rd_data_bits_9_9(load_io_wgt_rd_data_bits_9_9),
    .io_wgt_rd_data_bits_9_10(load_io_wgt_rd_data_bits_9_10),
    .io_wgt_rd_data_bits_9_11(load_io_wgt_rd_data_bits_9_11),
    .io_wgt_rd_data_bits_9_12(load_io_wgt_rd_data_bits_9_12),
    .io_wgt_rd_data_bits_9_13(load_io_wgt_rd_data_bits_9_13),
    .io_wgt_rd_data_bits_9_14(load_io_wgt_rd_data_bits_9_14),
    .io_wgt_rd_data_bits_9_15(load_io_wgt_rd_data_bits_9_15),
    .io_wgt_rd_data_bits_10_0(load_io_wgt_rd_data_bits_10_0),
    .io_wgt_rd_data_bits_10_1(load_io_wgt_rd_data_bits_10_1),
    .io_wgt_rd_data_bits_10_2(load_io_wgt_rd_data_bits_10_2),
    .io_wgt_rd_data_bits_10_3(load_io_wgt_rd_data_bits_10_3),
    .io_wgt_rd_data_bits_10_4(load_io_wgt_rd_data_bits_10_4),
    .io_wgt_rd_data_bits_10_5(load_io_wgt_rd_data_bits_10_5),
    .io_wgt_rd_data_bits_10_6(load_io_wgt_rd_data_bits_10_6),
    .io_wgt_rd_data_bits_10_7(load_io_wgt_rd_data_bits_10_7),
    .io_wgt_rd_data_bits_10_8(load_io_wgt_rd_data_bits_10_8),
    .io_wgt_rd_data_bits_10_9(load_io_wgt_rd_data_bits_10_9),
    .io_wgt_rd_data_bits_10_10(load_io_wgt_rd_data_bits_10_10),
    .io_wgt_rd_data_bits_10_11(load_io_wgt_rd_data_bits_10_11),
    .io_wgt_rd_data_bits_10_12(load_io_wgt_rd_data_bits_10_12),
    .io_wgt_rd_data_bits_10_13(load_io_wgt_rd_data_bits_10_13),
    .io_wgt_rd_data_bits_10_14(load_io_wgt_rd_data_bits_10_14),
    .io_wgt_rd_data_bits_10_15(load_io_wgt_rd_data_bits_10_15),
    .io_wgt_rd_data_bits_11_0(load_io_wgt_rd_data_bits_11_0),
    .io_wgt_rd_data_bits_11_1(load_io_wgt_rd_data_bits_11_1),
    .io_wgt_rd_data_bits_11_2(load_io_wgt_rd_data_bits_11_2),
    .io_wgt_rd_data_bits_11_3(load_io_wgt_rd_data_bits_11_3),
    .io_wgt_rd_data_bits_11_4(load_io_wgt_rd_data_bits_11_4),
    .io_wgt_rd_data_bits_11_5(load_io_wgt_rd_data_bits_11_5),
    .io_wgt_rd_data_bits_11_6(load_io_wgt_rd_data_bits_11_6),
    .io_wgt_rd_data_bits_11_7(load_io_wgt_rd_data_bits_11_7),
    .io_wgt_rd_data_bits_11_8(load_io_wgt_rd_data_bits_11_8),
    .io_wgt_rd_data_bits_11_9(load_io_wgt_rd_data_bits_11_9),
    .io_wgt_rd_data_bits_11_10(load_io_wgt_rd_data_bits_11_10),
    .io_wgt_rd_data_bits_11_11(load_io_wgt_rd_data_bits_11_11),
    .io_wgt_rd_data_bits_11_12(load_io_wgt_rd_data_bits_11_12),
    .io_wgt_rd_data_bits_11_13(load_io_wgt_rd_data_bits_11_13),
    .io_wgt_rd_data_bits_11_14(load_io_wgt_rd_data_bits_11_14),
    .io_wgt_rd_data_bits_11_15(load_io_wgt_rd_data_bits_11_15),
    .io_wgt_rd_data_bits_12_0(load_io_wgt_rd_data_bits_12_0),
    .io_wgt_rd_data_bits_12_1(load_io_wgt_rd_data_bits_12_1),
    .io_wgt_rd_data_bits_12_2(load_io_wgt_rd_data_bits_12_2),
    .io_wgt_rd_data_bits_12_3(load_io_wgt_rd_data_bits_12_3),
    .io_wgt_rd_data_bits_12_4(load_io_wgt_rd_data_bits_12_4),
    .io_wgt_rd_data_bits_12_5(load_io_wgt_rd_data_bits_12_5),
    .io_wgt_rd_data_bits_12_6(load_io_wgt_rd_data_bits_12_6),
    .io_wgt_rd_data_bits_12_7(load_io_wgt_rd_data_bits_12_7),
    .io_wgt_rd_data_bits_12_8(load_io_wgt_rd_data_bits_12_8),
    .io_wgt_rd_data_bits_12_9(load_io_wgt_rd_data_bits_12_9),
    .io_wgt_rd_data_bits_12_10(load_io_wgt_rd_data_bits_12_10),
    .io_wgt_rd_data_bits_12_11(load_io_wgt_rd_data_bits_12_11),
    .io_wgt_rd_data_bits_12_12(load_io_wgt_rd_data_bits_12_12),
    .io_wgt_rd_data_bits_12_13(load_io_wgt_rd_data_bits_12_13),
    .io_wgt_rd_data_bits_12_14(load_io_wgt_rd_data_bits_12_14),
    .io_wgt_rd_data_bits_12_15(load_io_wgt_rd_data_bits_12_15),
    .io_wgt_rd_data_bits_13_0(load_io_wgt_rd_data_bits_13_0),
    .io_wgt_rd_data_bits_13_1(load_io_wgt_rd_data_bits_13_1),
    .io_wgt_rd_data_bits_13_2(load_io_wgt_rd_data_bits_13_2),
    .io_wgt_rd_data_bits_13_3(load_io_wgt_rd_data_bits_13_3),
    .io_wgt_rd_data_bits_13_4(load_io_wgt_rd_data_bits_13_4),
    .io_wgt_rd_data_bits_13_5(load_io_wgt_rd_data_bits_13_5),
    .io_wgt_rd_data_bits_13_6(load_io_wgt_rd_data_bits_13_6),
    .io_wgt_rd_data_bits_13_7(load_io_wgt_rd_data_bits_13_7),
    .io_wgt_rd_data_bits_13_8(load_io_wgt_rd_data_bits_13_8),
    .io_wgt_rd_data_bits_13_9(load_io_wgt_rd_data_bits_13_9),
    .io_wgt_rd_data_bits_13_10(load_io_wgt_rd_data_bits_13_10),
    .io_wgt_rd_data_bits_13_11(load_io_wgt_rd_data_bits_13_11),
    .io_wgt_rd_data_bits_13_12(load_io_wgt_rd_data_bits_13_12),
    .io_wgt_rd_data_bits_13_13(load_io_wgt_rd_data_bits_13_13),
    .io_wgt_rd_data_bits_13_14(load_io_wgt_rd_data_bits_13_14),
    .io_wgt_rd_data_bits_13_15(load_io_wgt_rd_data_bits_13_15),
    .io_wgt_rd_data_bits_14_0(load_io_wgt_rd_data_bits_14_0),
    .io_wgt_rd_data_bits_14_1(load_io_wgt_rd_data_bits_14_1),
    .io_wgt_rd_data_bits_14_2(load_io_wgt_rd_data_bits_14_2),
    .io_wgt_rd_data_bits_14_3(load_io_wgt_rd_data_bits_14_3),
    .io_wgt_rd_data_bits_14_4(load_io_wgt_rd_data_bits_14_4),
    .io_wgt_rd_data_bits_14_5(load_io_wgt_rd_data_bits_14_5),
    .io_wgt_rd_data_bits_14_6(load_io_wgt_rd_data_bits_14_6),
    .io_wgt_rd_data_bits_14_7(load_io_wgt_rd_data_bits_14_7),
    .io_wgt_rd_data_bits_14_8(load_io_wgt_rd_data_bits_14_8),
    .io_wgt_rd_data_bits_14_9(load_io_wgt_rd_data_bits_14_9),
    .io_wgt_rd_data_bits_14_10(load_io_wgt_rd_data_bits_14_10),
    .io_wgt_rd_data_bits_14_11(load_io_wgt_rd_data_bits_14_11),
    .io_wgt_rd_data_bits_14_12(load_io_wgt_rd_data_bits_14_12),
    .io_wgt_rd_data_bits_14_13(load_io_wgt_rd_data_bits_14_13),
    .io_wgt_rd_data_bits_14_14(load_io_wgt_rd_data_bits_14_14),
    .io_wgt_rd_data_bits_14_15(load_io_wgt_rd_data_bits_14_15),
    .io_wgt_rd_data_bits_15_0(load_io_wgt_rd_data_bits_15_0),
    .io_wgt_rd_data_bits_15_1(load_io_wgt_rd_data_bits_15_1),
    .io_wgt_rd_data_bits_15_2(load_io_wgt_rd_data_bits_15_2),
    .io_wgt_rd_data_bits_15_3(load_io_wgt_rd_data_bits_15_3),
    .io_wgt_rd_data_bits_15_4(load_io_wgt_rd_data_bits_15_4),
    .io_wgt_rd_data_bits_15_5(load_io_wgt_rd_data_bits_15_5),
    .io_wgt_rd_data_bits_15_6(load_io_wgt_rd_data_bits_15_6),
    .io_wgt_rd_data_bits_15_7(load_io_wgt_rd_data_bits_15_7),
    .io_wgt_rd_data_bits_15_8(load_io_wgt_rd_data_bits_15_8),
    .io_wgt_rd_data_bits_15_9(load_io_wgt_rd_data_bits_15_9),
    .io_wgt_rd_data_bits_15_10(load_io_wgt_rd_data_bits_15_10),
    .io_wgt_rd_data_bits_15_11(load_io_wgt_rd_data_bits_15_11),
    .io_wgt_rd_data_bits_15_12(load_io_wgt_rd_data_bits_15_12),
    .io_wgt_rd_data_bits_15_13(load_io_wgt_rd_data_bits_15_13),
    .io_wgt_rd_data_bits_15_14(load_io_wgt_rd_data_bits_15_14),
    .io_wgt_rd_data_bits_15_15(load_io_wgt_rd_data_bits_15_15)
  );
  Compute compute ( // @[Core.scala 68:23:@24758.4]
    .clock(compute_clock),
    .reset(compute_reset),
    .io_i_post_0(compute_io_i_post_0),
    .io_i_post_1(compute_io_i_post_1),
    .io_o_post_0(compute_io_o_post_0),
    .io_o_post_1(compute_io_o_post_1),
    .io_inst_ready(compute_io_inst_ready),
    .io_inst_valid(compute_io_inst_valid),
    .io_inst_bits(compute_io_inst_bits),
    .io_uop_baddr(compute_io_uop_baddr),
    .io_acc_baddr(compute_io_acc_baddr),
    .io_vme_rd_0_cmd_ready(compute_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(compute_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(compute_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(compute_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(compute_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(compute_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits(compute_io_vme_rd_0_data_bits),
    .io_vme_rd_1_cmd_ready(compute_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(compute_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(compute_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(compute_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_data_ready(compute_io_vme_rd_1_data_ready),
    .io_vme_rd_1_data_valid(compute_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits(compute_io_vme_rd_1_data_bits),
    .io_inp_rd_idx_valid(compute_io_inp_rd_idx_valid),
    .io_inp_rd_idx_bits(compute_io_inp_rd_idx_bits),
    .io_inp_rd_data_valid(compute_io_inp_rd_data_valid),
    .io_inp_rd_data_bits_0_0(compute_io_inp_rd_data_bits_0_0),
    .io_inp_rd_data_bits_0_1(compute_io_inp_rd_data_bits_0_1),
    .io_inp_rd_data_bits_0_2(compute_io_inp_rd_data_bits_0_2),
    .io_inp_rd_data_bits_0_3(compute_io_inp_rd_data_bits_0_3),
    .io_inp_rd_data_bits_0_4(compute_io_inp_rd_data_bits_0_4),
    .io_inp_rd_data_bits_0_5(compute_io_inp_rd_data_bits_0_5),
    .io_inp_rd_data_bits_0_6(compute_io_inp_rd_data_bits_0_6),
    .io_inp_rd_data_bits_0_7(compute_io_inp_rd_data_bits_0_7),
    .io_inp_rd_data_bits_0_8(compute_io_inp_rd_data_bits_0_8),
    .io_inp_rd_data_bits_0_9(compute_io_inp_rd_data_bits_0_9),
    .io_inp_rd_data_bits_0_10(compute_io_inp_rd_data_bits_0_10),
    .io_inp_rd_data_bits_0_11(compute_io_inp_rd_data_bits_0_11),
    .io_inp_rd_data_bits_0_12(compute_io_inp_rd_data_bits_0_12),
    .io_inp_rd_data_bits_0_13(compute_io_inp_rd_data_bits_0_13),
    .io_inp_rd_data_bits_0_14(compute_io_inp_rd_data_bits_0_14),
    .io_inp_rd_data_bits_0_15(compute_io_inp_rd_data_bits_0_15),
    .io_wgt_rd_idx_valid(compute_io_wgt_rd_idx_valid),
    .io_wgt_rd_idx_bits(compute_io_wgt_rd_idx_bits),
    .io_wgt_rd_data_valid(compute_io_wgt_rd_data_valid),
    .io_wgt_rd_data_bits_0_0(compute_io_wgt_rd_data_bits_0_0),
    .io_wgt_rd_data_bits_0_1(compute_io_wgt_rd_data_bits_0_1),
    .io_wgt_rd_data_bits_0_2(compute_io_wgt_rd_data_bits_0_2),
    .io_wgt_rd_data_bits_0_3(compute_io_wgt_rd_data_bits_0_3),
    .io_wgt_rd_data_bits_0_4(compute_io_wgt_rd_data_bits_0_4),
    .io_wgt_rd_data_bits_0_5(compute_io_wgt_rd_data_bits_0_5),
    .io_wgt_rd_data_bits_0_6(compute_io_wgt_rd_data_bits_0_6),
    .io_wgt_rd_data_bits_0_7(compute_io_wgt_rd_data_bits_0_7),
    .io_wgt_rd_data_bits_0_8(compute_io_wgt_rd_data_bits_0_8),
    .io_wgt_rd_data_bits_0_9(compute_io_wgt_rd_data_bits_0_9),
    .io_wgt_rd_data_bits_0_10(compute_io_wgt_rd_data_bits_0_10),
    .io_wgt_rd_data_bits_0_11(compute_io_wgt_rd_data_bits_0_11),
    .io_wgt_rd_data_bits_0_12(compute_io_wgt_rd_data_bits_0_12),
    .io_wgt_rd_data_bits_0_13(compute_io_wgt_rd_data_bits_0_13),
    .io_wgt_rd_data_bits_0_14(compute_io_wgt_rd_data_bits_0_14),
    .io_wgt_rd_data_bits_0_15(compute_io_wgt_rd_data_bits_0_15),
    .io_wgt_rd_data_bits_1_0(compute_io_wgt_rd_data_bits_1_0),
    .io_wgt_rd_data_bits_1_1(compute_io_wgt_rd_data_bits_1_1),
    .io_wgt_rd_data_bits_1_2(compute_io_wgt_rd_data_bits_1_2),
    .io_wgt_rd_data_bits_1_3(compute_io_wgt_rd_data_bits_1_3),
    .io_wgt_rd_data_bits_1_4(compute_io_wgt_rd_data_bits_1_4),
    .io_wgt_rd_data_bits_1_5(compute_io_wgt_rd_data_bits_1_5),
    .io_wgt_rd_data_bits_1_6(compute_io_wgt_rd_data_bits_1_6),
    .io_wgt_rd_data_bits_1_7(compute_io_wgt_rd_data_bits_1_7),
    .io_wgt_rd_data_bits_1_8(compute_io_wgt_rd_data_bits_1_8),
    .io_wgt_rd_data_bits_1_9(compute_io_wgt_rd_data_bits_1_9),
    .io_wgt_rd_data_bits_1_10(compute_io_wgt_rd_data_bits_1_10),
    .io_wgt_rd_data_bits_1_11(compute_io_wgt_rd_data_bits_1_11),
    .io_wgt_rd_data_bits_1_12(compute_io_wgt_rd_data_bits_1_12),
    .io_wgt_rd_data_bits_1_13(compute_io_wgt_rd_data_bits_1_13),
    .io_wgt_rd_data_bits_1_14(compute_io_wgt_rd_data_bits_1_14),
    .io_wgt_rd_data_bits_1_15(compute_io_wgt_rd_data_bits_1_15),
    .io_wgt_rd_data_bits_2_0(compute_io_wgt_rd_data_bits_2_0),
    .io_wgt_rd_data_bits_2_1(compute_io_wgt_rd_data_bits_2_1),
    .io_wgt_rd_data_bits_2_2(compute_io_wgt_rd_data_bits_2_2),
    .io_wgt_rd_data_bits_2_3(compute_io_wgt_rd_data_bits_2_3),
    .io_wgt_rd_data_bits_2_4(compute_io_wgt_rd_data_bits_2_4),
    .io_wgt_rd_data_bits_2_5(compute_io_wgt_rd_data_bits_2_5),
    .io_wgt_rd_data_bits_2_6(compute_io_wgt_rd_data_bits_2_6),
    .io_wgt_rd_data_bits_2_7(compute_io_wgt_rd_data_bits_2_7),
    .io_wgt_rd_data_bits_2_8(compute_io_wgt_rd_data_bits_2_8),
    .io_wgt_rd_data_bits_2_9(compute_io_wgt_rd_data_bits_2_9),
    .io_wgt_rd_data_bits_2_10(compute_io_wgt_rd_data_bits_2_10),
    .io_wgt_rd_data_bits_2_11(compute_io_wgt_rd_data_bits_2_11),
    .io_wgt_rd_data_bits_2_12(compute_io_wgt_rd_data_bits_2_12),
    .io_wgt_rd_data_bits_2_13(compute_io_wgt_rd_data_bits_2_13),
    .io_wgt_rd_data_bits_2_14(compute_io_wgt_rd_data_bits_2_14),
    .io_wgt_rd_data_bits_2_15(compute_io_wgt_rd_data_bits_2_15),
    .io_wgt_rd_data_bits_3_0(compute_io_wgt_rd_data_bits_3_0),
    .io_wgt_rd_data_bits_3_1(compute_io_wgt_rd_data_bits_3_1),
    .io_wgt_rd_data_bits_3_2(compute_io_wgt_rd_data_bits_3_2),
    .io_wgt_rd_data_bits_3_3(compute_io_wgt_rd_data_bits_3_3),
    .io_wgt_rd_data_bits_3_4(compute_io_wgt_rd_data_bits_3_4),
    .io_wgt_rd_data_bits_3_5(compute_io_wgt_rd_data_bits_3_5),
    .io_wgt_rd_data_bits_3_6(compute_io_wgt_rd_data_bits_3_6),
    .io_wgt_rd_data_bits_3_7(compute_io_wgt_rd_data_bits_3_7),
    .io_wgt_rd_data_bits_3_8(compute_io_wgt_rd_data_bits_3_8),
    .io_wgt_rd_data_bits_3_9(compute_io_wgt_rd_data_bits_3_9),
    .io_wgt_rd_data_bits_3_10(compute_io_wgt_rd_data_bits_3_10),
    .io_wgt_rd_data_bits_3_11(compute_io_wgt_rd_data_bits_3_11),
    .io_wgt_rd_data_bits_3_12(compute_io_wgt_rd_data_bits_3_12),
    .io_wgt_rd_data_bits_3_13(compute_io_wgt_rd_data_bits_3_13),
    .io_wgt_rd_data_bits_3_14(compute_io_wgt_rd_data_bits_3_14),
    .io_wgt_rd_data_bits_3_15(compute_io_wgt_rd_data_bits_3_15),
    .io_wgt_rd_data_bits_4_0(compute_io_wgt_rd_data_bits_4_0),
    .io_wgt_rd_data_bits_4_1(compute_io_wgt_rd_data_bits_4_1),
    .io_wgt_rd_data_bits_4_2(compute_io_wgt_rd_data_bits_4_2),
    .io_wgt_rd_data_bits_4_3(compute_io_wgt_rd_data_bits_4_3),
    .io_wgt_rd_data_bits_4_4(compute_io_wgt_rd_data_bits_4_4),
    .io_wgt_rd_data_bits_4_5(compute_io_wgt_rd_data_bits_4_5),
    .io_wgt_rd_data_bits_4_6(compute_io_wgt_rd_data_bits_4_6),
    .io_wgt_rd_data_bits_4_7(compute_io_wgt_rd_data_bits_4_7),
    .io_wgt_rd_data_bits_4_8(compute_io_wgt_rd_data_bits_4_8),
    .io_wgt_rd_data_bits_4_9(compute_io_wgt_rd_data_bits_4_9),
    .io_wgt_rd_data_bits_4_10(compute_io_wgt_rd_data_bits_4_10),
    .io_wgt_rd_data_bits_4_11(compute_io_wgt_rd_data_bits_4_11),
    .io_wgt_rd_data_bits_4_12(compute_io_wgt_rd_data_bits_4_12),
    .io_wgt_rd_data_bits_4_13(compute_io_wgt_rd_data_bits_4_13),
    .io_wgt_rd_data_bits_4_14(compute_io_wgt_rd_data_bits_4_14),
    .io_wgt_rd_data_bits_4_15(compute_io_wgt_rd_data_bits_4_15),
    .io_wgt_rd_data_bits_5_0(compute_io_wgt_rd_data_bits_5_0),
    .io_wgt_rd_data_bits_5_1(compute_io_wgt_rd_data_bits_5_1),
    .io_wgt_rd_data_bits_5_2(compute_io_wgt_rd_data_bits_5_2),
    .io_wgt_rd_data_bits_5_3(compute_io_wgt_rd_data_bits_5_3),
    .io_wgt_rd_data_bits_5_4(compute_io_wgt_rd_data_bits_5_4),
    .io_wgt_rd_data_bits_5_5(compute_io_wgt_rd_data_bits_5_5),
    .io_wgt_rd_data_bits_5_6(compute_io_wgt_rd_data_bits_5_6),
    .io_wgt_rd_data_bits_5_7(compute_io_wgt_rd_data_bits_5_7),
    .io_wgt_rd_data_bits_5_8(compute_io_wgt_rd_data_bits_5_8),
    .io_wgt_rd_data_bits_5_9(compute_io_wgt_rd_data_bits_5_9),
    .io_wgt_rd_data_bits_5_10(compute_io_wgt_rd_data_bits_5_10),
    .io_wgt_rd_data_bits_5_11(compute_io_wgt_rd_data_bits_5_11),
    .io_wgt_rd_data_bits_5_12(compute_io_wgt_rd_data_bits_5_12),
    .io_wgt_rd_data_bits_5_13(compute_io_wgt_rd_data_bits_5_13),
    .io_wgt_rd_data_bits_5_14(compute_io_wgt_rd_data_bits_5_14),
    .io_wgt_rd_data_bits_5_15(compute_io_wgt_rd_data_bits_5_15),
    .io_wgt_rd_data_bits_6_0(compute_io_wgt_rd_data_bits_6_0),
    .io_wgt_rd_data_bits_6_1(compute_io_wgt_rd_data_bits_6_1),
    .io_wgt_rd_data_bits_6_2(compute_io_wgt_rd_data_bits_6_2),
    .io_wgt_rd_data_bits_6_3(compute_io_wgt_rd_data_bits_6_3),
    .io_wgt_rd_data_bits_6_4(compute_io_wgt_rd_data_bits_6_4),
    .io_wgt_rd_data_bits_6_5(compute_io_wgt_rd_data_bits_6_5),
    .io_wgt_rd_data_bits_6_6(compute_io_wgt_rd_data_bits_6_6),
    .io_wgt_rd_data_bits_6_7(compute_io_wgt_rd_data_bits_6_7),
    .io_wgt_rd_data_bits_6_8(compute_io_wgt_rd_data_bits_6_8),
    .io_wgt_rd_data_bits_6_9(compute_io_wgt_rd_data_bits_6_9),
    .io_wgt_rd_data_bits_6_10(compute_io_wgt_rd_data_bits_6_10),
    .io_wgt_rd_data_bits_6_11(compute_io_wgt_rd_data_bits_6_11),
    .io_wgt_rd_data_bits_6_12(compute_io_wgt_rd_data_bits_6_12),
    .io_wgt_rd_data_bits_6_13(compute_io_wgt_rd_data_bits_6_13),
    .io_wgt_rd_data_bits_6_14(compute_io_wgt_rd_data_bits_6_14),
    .io_wgt_rd_data_bits_6_15(compute_io_wgt_rd_data_bits_6_15),
    .io_wgt_rd_data_bits_7_0(compute_io_wgt_rd_data_bits_7_0),
    .io_wgt_rd_data_bits_7_1(compute_io_wgt_rd_data_bits_7_1),
    .io_wgt_rd_data_bits_7_2(compute_io_wgt_rd_data_bits_7_2),
    .io_wgt_rd_data_bits_7_3(compute_io_wgt_rd_data_bits_7_3),
    .io_wgt_rd_data_bits_7_4(compute_io_wgt_rd_data_bits_7_4),
    .io_wgt_rd_data_bits_7_5(compute_io_wgt_rd_data_bits_7_5),
    .io_wgt_rd_data_bits_7_6(compute_io_wgt_rd_data_bits_7_6),
    .io_wgt_rd_data_bits_7_7(compute_io_wgt_rd_data_bits_7_7),
    .io_wgt_rd_data_bits_7_8(compute_io_wgt_rd_data_bits_7_8),
    .io_wgt_rd_data_bits_7_9(compute_io_wgt_rd_data_bits_7_9),
    .io_wgt_rd_data_bits_7_10(compute_io_wgt_rd_data_bits_7_10),
    .io_wgt_rd_data_bits_7_11(compute_io_wgt_rd_data_bits_7_11),
    .io_wgt_rd_data_bits_7_12(compute_io_wgt_rd_data_bits_7_12),
    .io_wgt_rd_data_bits_7_13(compute_io_wgt_rd_data_bits_7_13),
    .io_wgt_rd_data_bits_7_14(compute_io_wgt_rd_data_bits_7_14),
    .io_wgt_rd_data_bits_7_15(compute_io_wgt_rd_data_bits_7_15),
    .io_wgt_rd_data_bits_8_0(compute_io_wgt_rd_data_bits_8_0),
    .io_wgt_rd_data_bits_8_1(compute_io_wgt_rd_data_bits_8_1),
    .io_wgt_rd_data_bits_8_2(compute_io_wgt_rd_data_bits_8_2),
    .io_wgt_rd_data_bits_8_3(compute_io_wgt_rd_data_bits_8_3),
    .io_wgt_rd_data_bits_8_4(compute_io_wgt_rd_data_bits_8_4),
    .io_wgt_rd_data_bits_8_5(compute_io_wgt_rd_data_bits_8_5),
    .io_wgt_rd_data_bits_8_6(compute_io_wgt_rd_data_bits_8_6),
    .io_wgt_rd_data_bits_8_7(compute_io_wgt_rd_data_bits_8_7),
    .io_wgt_rd_data_bits_8_8(compute_io_wgt_rd_data_bits_8_8),
    .io_wgt_rd_data_bits_8_9(compute_io_wgt_rd_data_bits_8_9),
    .io_wgt_rd_data_bits_8_10(compute_io_wgt_rd_data_bits_8_10),
    .io_wgt_rd_data_bits_8_11(compute_io_wgt_rd_data_bits_8_11),
    .io_wgt_rd_data_bits_8_12(compute_io_wgt_rd_data_bits_8_12),
    .io_wgt_rd_data_bits_8_13(compute_io_wgt_rd_data_bits_8_13),
    .io_wgt_rd_data_bits_8_14(compute_io_wgt_rd_data_bits_8_14),
    .io_wgt_rd_data_bits_8_15(compute_io_wgt_rd_data_bits_8_15),
    .io_wgt_rd_data_bits_9_0(compute_io_wgt_rd_data_bits_9_0),
    .io_wgt_rd_data_bits_9_1(compute_io_wgt_rd_data_bits_9_1),
    .io_wgt_rd_data_bits_9_2(compute_io_wgt_rd_data_bits_9_2),
    .io_wgt_rd_data_bits_9_3(compute_io_wgt_rd_data_bits_9_3),
    .io_wgt_rd_data_bits_9_4(compute_io_wgt_rd_data_bits_9_4),
    .io_wgt_rd_data_bits_9_5(compute_io_wgt_rd_data_bits_9_5),
    .io_wgt_rd_data_bits_9_6(compute_io_wgt_rd_data_bits_9_6),
    .io_wgt_rd_data_bits_9_7(compute_io_wgt_rd_data_bits_9_7),
    .io_wgt_rd_data_bits_9_8(compute_io_wgt_rd_data_bits_9_8),
    .io_wgt_rd_data_bits_9_9(compute_io_wgt_rd_data_bits_9_9),
    .io_wgt_rd_data_bits_9_10(compute_io_wgt_rd_data_bits_9_10),
    .io_wgt_rd_data_bits_9_11(compute_io_wgt_rd_data_bits_9_11),
    .io_wgt_rd_data_bits_9_12(compute_io_wgt_rd_data_bits_9_12),
    .io_wgt_rd_data_bits_9_13(compute_io_wgt_rd_data_bits_9_13),
    .io_wgt_rd_data_bits_9_14(compute_io_wgt_rd_data_bits_9_14),
    .io_wgt_rd_data_bits_9_15(compute_io_wgt_rd_data_bits_9_15),
    .io_wgt_rd_data_bits_10_0(compute_io_wgt_rd_data_bits_10_0),
    .io_wgt_rd_data_bits_10_1(compute_io_wgt_rd_data_bits_10_1),
    .io_wgt_rd_data_bits_10_2(compute_io_wgt_rd_data_bits_10_2),
    .io_wgt_rd_data_bits_10_3(compute_io_wgt_rd_data_bits_10_3),
    .io_wgt_rd_data_bits_10_4(compute_io_wgt_rd_data_bits_10_4),
    .io_wgt_rd_data_bits_10_5(compute_io_wgt_rd_data_bits_10_5),
    .io_wgt_rd_data_bits_10_6(compute_io_wgt_rd_data_bits_10_6),
    .io_wgt_rd_data_bits_10_7(compute_io_wgt_rd_data_bits_10_7),
    .io_wgt_rd_data_bits_10_8(compute_io_wgt_rd_data_bits_10_8),
    .io_wgt_rd_data_bits_10_9(compute_io_wgt_rd_data_bits_10_9),
    .io_wgt_rd_data_bits_10_10(compute_io_wgt_rd_data_bits_10_10),
    .io_wgt_rd_data_bits_10_11(compute_io_wgt_rd_data_bits_10_11),
    .io_wgt_rd_data_bits_10_12(compute_io_wgt_rd_data_bits_10_12),
    .io_wgt_rd_data_bits_10_13(compute_io_wgt_rd_data_bits_10_13),
    .io_wgt_rd_data_bits_10_14(compute_io_wgt_rd_data_bits_10_14),
    .io_wgt_rd_data_bits_10_15(compute_io_wgt_rd_data_bits_10_15),
    .io_wgt_rd_data_bits_11_0(compute_io_wgt_rd_data_bits_11_0),
    .io_wgt_rd_data_bits_11_1(compute_io_wgt_rd_data_bits_11_1),
    .io_wgt_rd_data_bits_11_2(compute_io_wgt_rd_data_bits_11_2),
    .io_wgt_rd_data_bits_11_3(compute_io_wgt_rd_data_bits_11_3),
    .io_wgt_rd_data_bits_11_4(compute_io_wgt_rd_data_bits_11_4),
    .io_wgt_rd_data_bits_11_5(compute_io_wgt_rd_data_bits_11_5),
    .io_wgt_rd_data_bits_11_6(compute_io_wgt_rd_data_bits_11_6),
    .io_wgt_rd_data_bits_11_7(compute_io_wgt_rd_data_bits_11_7),
    .io_wgt_rd_data_bits_11_8(compute_io_wgt_rd_data_bits_11_8),
    .io_wgt_rd_data_bits_11_9(compute_io_wgt_rd_data_bits_11_9),
    .io_wgt_rd_data_bits_11_10(compute_io_wgt_rd_data_bits_11_10),
    .io_wgt_rd_data_bits_11_11(compute_io_wgt_rd_data_bits_11_11),
    .io_wgt_rd_data_bits_11_12(compute_io_wgt_rd_data_bits_11_12),
    .io_wgt_rd_data_bits_11_13(compute_io_wgt_rd_data_bits_11_13),
    .io_wgt_rd_data_bits_11_14(compute_io_wgt_rd_data_bits_11_14),
    .io_wgt_rd_data_bits_11_15(compute_io_wgt_rd_data_bits_11_15),
    .io_wgt_rd_data_bits_12_0(compute_io_wgt_rd_data_bits_12_0),
    .io_wgt_rd_data_bits_12_1(compute_io_wgt_rd_data_bits_12_1),
    .io_wgt_rd_data_bits_12_2(compute_io_wgt_rd_data_bits_12_2),
    .io_wgt_rd_data_bits_12_3(compute_io_wgt_rd_data_bits_12_3),
    .io_wgt_rd_data_bits_12_4(compute_io_wgt_rd_data_bits_12_4),
    .io_wgt_rd_data_bits_12_5(compute_io_wgt_rd_data_bits_12_5),
    .io_wgt_rd_data_bits_12_6(compute_io_wgt_rd_data_bits_12_6),
    .io_wgt_rd_data_bits_12_7(compute_io_wgt_rd_data_bits_12_7),
    .io_wgt_rd_data_bits_12_8(compute_io_wgt_rd_data_bits_12_8),
    .io_wgt_rd_data_bits_12_9(compute_io_wgt_rd_data_bits_12_9),
    .io_wgt_rd_data_bits_12_10(compute_io_wgt_rd_data_bits_12_10),
    .io_wgt_rd_data_bits_12_11(compute_io_wgt_rd_data_bits_12_11),
    .io_wgt_rd_data_bits_12_12(compute_io_wgt_rd_data_bits_12_12),
    .io_wgt_rd_data_bits_12_13(compute_io_wgt_rd_data_bits_12_13),
    .io_wgt_rd_data_bits_12_14(compute_io_wgt_rd_data_bits_12_14),
    .io_wgt_rd_data_bits_12_15(compute_io_wgt_rd_data_bits_12_15),
    .io_wgt_rd_data_bits_13_0(compute_io_wgt_rd_data_bits_13_0),
    .io_wgt_rd_data_bits_13_1(compute_io_wgt_rd_data_bits_13_1),
    .io_wgt_rd_data_bits_13_2(compute_io_wgt_rd_data_bits_13_2),
    .io_wgt_rd_data_bits_13_3(compute_io_wgt_rd_data_bits_13_3),
    .io_wgt_rd_data_bits_13_4(compute_io_wgt_rd_data_bits_13_4),
    .io_wgt_rd_data_bits_13_5(compute_io_wgt_rd_data_bits_13_5),
    .io_wgt_rd_data_bits_13_6(compute_io_wgt_rd_data_bits_13_6),
    .io_wgt_rd_data_bits_13_7(compute_io_wgt_rd_data_bits_13_7),
    .io_wgt_rd_data_bits_13_8(compute_io_wgt_rd_data_bits_13_8),
    .io_wgt_rd_data_bits_13_9(compute_io_wgt_rd_data_bits_13_9),
    .io_wgt_rd_data_bits_13_10(compute_io_wgt_rd_data_bits_13_10),
    .io_wgt_rd_data_bits_13_11(compute_io_wgt_rd_data_bits_13_11),
    .io_wgt_rd_data_bits_13_12(compute_io_wgt_rd_data_bits_13_12),
    .io_wgt_rd_data_bits_13_13(compute_io_wgt_rd_data_bits_13_13),
    .io_wgt_rd_data_bits_13_14(compute_io_wgt_rd_data_bits_13_14),
    .io_wgt_rd_data_bits_13_15(compute_io_wgt_rd_data_bits_13_15),
    .io_wgt_rd_data_bits_14_0(compute_io_wgt_rd_data_bits_14_0),
    .io_wgt_rd_data_bits_14_1(compute_io_wgt_rd_data_bits_14_1),
    .io_wgt_rd_data_bits_14_2(compute_io_wgt_rd_data_bits_14_2),
    .io_wgt_rd_data_bits_14_3(compute_io_wgt_rd_data_bits_14_3),
    .io_wgt_rd_data_bits_14_4(compute_io_wgt_rd_data_bits_14_4),
    .io_wgt_rd_data_bits_14_5(compute_io_wgt_rd_data_bits_14_5),
    .io_wgt_rd_data_bits_14_6(compute_io_wgt_rd_data_bits_14_6),
    .io_wgt_rd_data_bits_14_7(compute_io_wgt_rd_data_bits_14_7),
    .io_wgt_rd_data_bits_14_8(compute_io_wgt_rd_data_bits_14_8),
    .io_wgt_rd_data_bits_14_9(compute_io_wgt_rd_data_bits_14_9),
    .io_wgt_rd_data_bits_14_10(compute_io_wgt_rd_data_bits_14_10),
    .io_wgt_rd_data_bits_14_11(compute_io_wgt_rd_data_bits_14_11),
    .io_wgt_rd_data_bits_14_12(compute_io_wgt_rd_data_bits_14_12),
    .io_wgt_rd_data_bits_14_13(compute_io_wgt_rd_data_bits_14_13),
    .io_wgt_rd_data_bits_14_14(compute_io_wgt_rd_data_bits_14_14),
    .io_wgt_rd_data_bits_14_15(compute_io_wgt_rd_data_bits_14_15),
    .io_wgt_rd_data_bits_15_0(compute_io_wgt_rd_data_bits_15_0),
    .io_wgt_rd_data_bits_15_1(compute_io_wgt_rd_data_bits_15_1),
    .io_wgt_rd_data_bits_15_2(compute_io_wgt_rd_data_bits_15_2),
    .io_wgt_rd_data_bits_15_3(compute_io_wgt_rd_data_bits_15_3),
    .io_wgt_rd_data_bits_15_4(compute_io_wgt_rd_data_bits_15_4),
    .io_wgt_rd_data_bits_15_5(compute_io_wgt_rd_data_bits_15_5),
    .io_wgt_rd_data_bits_15_6(compute_io_wgt_rd_data_bits_15_6),
    .io_wgt_rd_data_bits_15_7(compute_io_wgt_rd_data_bits_15_7),
    .io_wgt_rd_data_bits_15_8(compute_io_wgt_rd_data_bits_15_8),
    .io_wgt_rd_data_bits_15_9(compute_io_wgt_rd_data_bits_15_9),
    .io_wgt_rd_data_bits_15_10(compute_io_wgt_rd_data_bits_15_10),
    .io_wgt_rd_data_bits_15_11(compute_io_wgt_rd_data_bits_15_11),
    .io_wgt_rd_data_bits_15_12(compute_io_wgt_rd_data_bits_15_12),
    .io_wgt_rd_data_bits_15_13(compute_io_wgt_rd_data_bits_15_13),
    .io_wgt_rd_data_bits_15_14(compute_io_wgt_rd_data_bits_15_14),
    .io_wgt_rd_data_bits_15_15(compute_io_wgt_rd_data_bits_15_15),
    .io_out_wr_valid(compute_io_out_wr_valid),
    .io_out_wr_bits_idx(compute_io_out_wr_bits_idx),
    .io_out_wr_bits_data_0_0(compute_io_out_wr_bits_data_0_0),
    .io_out_wr_bits_data_0_1(compute_io_out_wr_bits_data_0_1),
    .io_out_wr_bits_data_0_2(compute_io_out_wr_bits_data_0_2),
    .io_out_wr_bits_data_0_3(compute_io_out_wr_bits_data_0_3),
    .io_out_wr_bits_data_0_4(compute_io_out_wr_bits_data_0_4),
    .io_out_wr_bits_data_0_5(compute_io_out_wr_bits_data_0_5),
    .io_out_wr_bits_data_0_6(compute_io_out_wr_bits_data_0_6),
    .io_out_wr_bits_data_0_7(compute_io_out_wr_bits_data_0_7),
    .io_out_wr_bits_data_0_8(compute_io_out_wr_bits_data_0_8),
    .io_out_wr_bits_data_0_9(compute_io_out_wr_bits_data_0_9),
    .io_out_wr_bits_data_0_10(compute_io_out_wr_bits_data_0_10),
    .io_out_wr_bits_data_0_11(compute_io_out_wr_bits_data_0_11),
    .io_out_wr_bits_data_0_12(compute_io_out_wr_bits_data_0_12),
    .io_out_wr_bits_data_0_13(compute_io_out_wr_bits_data_0_13),
    .io_out_wr_bits_data_0_14(compute_io_out_wr_bits_data_0_14),
    .io_out_wr_bits_data_0_15(compute_io_out_wr_bits_data_0_15),
    .io_finish(compute_io_finish),
    .io_acc_wr_event(compute_io_acc_wr_event)
  );
  Store store ( // @[Core.scala 69:21:@24761.4]
    .clock(store_clock),
    .reset(store_reset),
    .io_i_post(store_io_i_post),
    .io_o_post(store_io_o_post),
    .io_inst_ready(store_io_inst_ready),
    .io_inst_valid(store_io_inst_valid),
    .io_inst_bits(store_io_inst_bits),
    .io_out_baddr(store_io_out_baddr),
    .io_vme_wr_cmd_ready(store_io_vme_wr_cmd_ready),
    .io_vme_wr_cmd_valid(store_io_vme_wr_cmd_valid),
    .io_vme_wr_cmd_bits_addr(store_io_vme_wr_cmd_bits_addr),
    .io_vme_wr_cmd_bits_len(store_io_vme_wr_cmd_bits_len),
    .io_vme_wr_data_ready(store_io_vme_wr_data_ready),
    .io_vme_wr_data_valid(store_io_vme_wr_data_valid),
    .io_vme_wr_data_bits(store_io_vme_wr_data_bits),
    .io_vme_wr_ack(store_io_vme_wr_ack),
    .io_out_wr_valid(store_io_out_wr_valid),
    .io_out_wr_bits_idx(store_io_out_wr_bits_idx),
    .io_out_wr_bits_data_0_0(store_io_out_wr_bits_data_0_0),
    .io_out_wr_bits_data_0_1(store_io_out_wr_bits_data_0_1),
    .io_out_wr_bits_data_0_2(store_io_out_wr_bits_data_0_2),
    .io_out_wr_bits_data_0_3(store_io_out_wr_bits_data_0_3),
    .io_out_wr_bits_data_0_4(store_io_out_wr_bits_data_0_4),
    .io_out_wr_bits_data_0_5(store_io_out_wr_bits_data_0_5),
    .io_out_wr_bits_data_0_6(store_io_out_wr_bits_data_0_6),
    .io_out_wr_bits_data_0_7(store_io_out_wr_bits_data_0_7),
    .io_out_wr_bits_data_0_8(store_io_out_wr_bits_data_0_8),
    .io_out_wr_bits_data_0_9(store_io_out_wr_bits_data_0_9),
    .io_out_wr_bits_data_0_10(store_io_out_wr_bits_data_0_10),
    .io_out_wr_bits_data_0_11(store_io_out_wr_bits_data_0_11),
    .io_out_wr_bits_data_0_12(store_io_out_wr_bits_data_0_12),
    .io_out_wr_bits_data_0_13(store_io_out_wr_bits_data_0_13),
    .io_out_wr_bits_data_0_14(store_io_out_wr_bits_data_0_14),
    .io_out_wr_bits_data_0_15(store_io_out_wr_bits_data_0_15)
  );
  EventCounters ecounters ( // @[Core.scala 70:25:@24764.4]
    .clock(ecounters_clock),
    .reset(ecounters_reset),
    .io_launch(ecounters_io_launch),
    .io_finish(ecounters_io_finish),
    .io_ecnt_0_valid(ecounters_io_ecnt_0_valid),
    .io_ecnt_0_bits(ecounters_io_ecnt_0_bits),
    .io_ucnt_0_valid(ecounters_io_ucnt_0_valid),
    .io_ucnt_0_bits(ecounters_io_ucnt_0_bits),
    .io_acc_wr_event(ecounters_io_acc_wr_event)
  );
  assign io_vcr_finish = finish; // @[Core.scala 119:17:@25431.4]
  assign io_vcr_ecnt_0_valid = ecounters_io_ecnt_0_valid; // @[Core.scala 113:15:@25425.4]
  assign io_vcr_ecnt_0_bits = ecounters_io_ecnt_0_bits; // @[Core.scala 113:15:@25424.4]
  assign io_vcr_ucnt_0_valid = ecounters_io_ucnt_0_valid; // @[Core.scala 114:15:@25427.4]
  assign io_vcr_ucnt_0_bits = ecounters_io_ucnt_0_bits; // @[Core.scala 114:15:@25426.4]
  assign io_vme_rd_0_cmd_valid = fetch_io_vme_rd_cmd_valid; // @[Core.scala 73:16:@24772.4]
  assign io_vme_rd_0_cmd_bits_addr = fetch_io_vme_rd_cmd_bits_addr; // @[Core.scala 73:16:@24771.4]
  assign io_vme_rd_0_cmd_bits_len = fetch_io_vme_rd_cmd_bits_len; // @[Core.scala 73:16:@24770.4]
  assign io_vme_rd_0_data_ready = fetch_io_vme_rd_data_ready; // @[Core.scala 73:16:@24769.4]
  assign io_vme_rd_1_cmd_valid = compute_io_vme_rd_0_cmd_valid; // @[Core.scala 74:16:@24779.4]
  assign io_vme_rd_1_cmd_bits_addr = compute_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 74:16:@24778.4]
  assign io_vme_rd_1_cmd_bits_len = compute_io_vme_rd_0_cmd_bits_len; // @[Core.scala 74:16:@24777.4]
  assign io_vme_rd_1_data_ready = compute_io_vme_rd_0_data_ready; // @[Core.scala 74:16:@24776.4]
  assign io_vme_rd_2_cmd_valid = load_io_vme_rd_0_cmd_valid; // @[Core.scala 75:16:@24786.4]
  assign io_vme_rd_2_cmd_bits_addr = load_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 75:16:@24785.4]
  assign io_vme_rd_2_cmd_bits_len = load_io_vme_rd_0_cmd_bits_len; // @[Core.scala 75:16:@24784.4]
  assign io_vme_rd_2_data_ready = load_io_vme_rd_0_data_ready; // @[Core.scala 75:16:@24783.4]
  assign io_vme_rd_3_cmd_valid = load_io_vme_rd_1_cmd_valid; // @[Core.scala 76:16:@24793.4]
  assign io_vme_rd_3_cmd_bits_addr = load_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 76:16:@24792.4]
  assign io_vme_rd_3_cmd_bits_len = load_io_vme_rd_1_cmd_bits_len; // @[Core.scala 76:16:@24791.4]
  assign io_vme_rd_3_data_ready = load_io_vme_rd_1_data_ready; // @[Core.scala 76:16:@24790.4]
  assign io_vme_rd_4_cmd_valid = compute_io_vme_rd_1_cmd_valid; // @[Core.scala 77:16:@24800.4]
  assign io_vme_rd_4_cmd_bits_addr = compute_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 77:16:@24799.4]
  assign io_vme_rd_4_cmd_bits_len = compute_io_vme_rd_1_cmd_bits_len; // @[Core.scala 77:16:@24798.4]
  assign io_vme_rd_4_data_ready = compute_io_vme_rd_1_data_ready; // @[Core.scala 77:16:@24797.4]
  assign io_vme_wr_0_cmd_valid = store_io_vme_wr_cmd_valid; // @[Core.scala 78:16:@24808.4]
  assign io_vme_wr_0_cmd_bits_addr = store_io_vme_wr_cmd_bits_addr; // @[Core.scala 78:16:@24807.4]
  assign io_vme_wr_0_cmd_bits_len = store_io_vme_wr_cmd_bits_len; // @[Core.scala 78:16:@24806.4]
  assign io_vme_wr_0_data_valid = store_io_vme_wr_data_valid; // @[Core.scala 78:16:@24804.4]
  assign io_vme_wr_0_data_bits = store_io_vme_wr_data_bits; // @[Core.scala 78:16:@24803.4]
  assign fetch_clock = clock; // @[:@24753.4]
  assign fetch_reset = reset; // @[:@24754.4]
  assign fetch_io_launch = io_vcr_launch; // @[Core.scala 81:19:@24810.4]
  assign fetch_io_ins_baddr = io_vcr_ptrs_0; // @[Core.scala 82:22:@24811.4]
  assign fetch_io_ins_count = io_vcr_vals_0; // @[Core.scala 83:22:@24812.4]
  assign fetch_io_vme_rd_cmd_ready = io_vme_rd_0_cmd_ready; // @[Core.scala 73:16:@24773.4]
  assign fetch_io_vme_rd_data_valid = io_vme_rd_0_data_valid; // @[Core.scala 73:16:@24768.4]
  assign fetch_io_vme_rd_data_bits = io_vme_rd_0_data_bits; // @[Core.scala 73:16:@24767.4]
  assign fetch_io_inst_ld_ready = load_io_inst_ready; // @[Core.scala 87:16:@24816.4]
  assign fetch_io_inst_co_ready = compute_io_inst_ready; // @[Core.scala 96:19:@24823.4]
  assign fetch_io_inst_st_ready = store_io_inst_ready; // @[Core.scala 106:17:@25383.4]
  assign load_clock = clock; // @[:@24756.4]
  assign load_reset = reset; // @[:@24757.4]
  assign load_io_i_post = compute_io_o_post_0; // @[Core.scala 86:18:@24813.4]
  assign load_io_inst_valid = fetch_io_inst_ld_valid; // @[Core.scala 87:16:@24815.4]
  assign load_io_inst_bits = fetch_io_inst_ld_bits; // @[Core.scala 87:16:@24814.4]
  assign load_io_inp_baddr = io_vcr_ptrs_2; // @[Core.scala 88:21:@24817.4]
  assign load_io_wgt_baddr = io_vcr_ptrs_3; // @[Core.scala 89:21:@24818.4]
  assign load_io_vme_rd_0_cmd_ready = io_vme_rd_2_cmd_ready; // @[Core.scala 75:16:@24787.4]
  assign load_io_vme_rd_0_data_valid = io_vme_rd_2_data_valid; // @[Core.scala 75:16:@24782.4]
  assign load_io_vme_rd_0_data_bits = io_vme_rd_2_data_bits; // @[Core.scala 75:16:@24781.4]
  assign load_io_vme_rd_1_cmd_ready = io_vme_rd_3_cmd_ready; // @[Core.scala 76:16:@24794.4]
  assign load_io_vme_rd_1_data_valid = io_vme_rd_3_data_valid; // @[Core.scala 76:16:@24789.4]
  assign load_io_vme_rd_1_data_bits = io_vme_rd_3_data_bits; // @[Core.scala 76:16:@24788.4]
  assign load_io_inp_rd_idx_valid = compute_io_inp_rd_idx_valid; // @[Core.scala 99:18:@24862.4]
  assign load_io_inp_rd_idx_bits = compute_io_inp_rd_idx_bits; // @[Core.scala 99:18:@24861.4]
  assign load_io_wgt_rd_idx_valid = compute_io_wgt_rd_idx_valid; // @[Core.scala 100:18:@25379.4]
  assign load_io_wgt_rd_idx_bits = compute_io_wgt_rd_idx_bits; // @[Core.scala 100:18:@25378.4]
  assign compute_clock = clock; // @[:@24759.4]
  assign compute_reset = reset; // @[:@24760.4]
  assign compute_io_i_post_0 = load_io_o_post; // @[Core.scala 94:24:@24819.4]
  assign compute_io_i_post_1 = store_io_o_post; // @[Core.scala 95:24:@24820.4]
  assign compute_io_inst_valid = fetch_io_inst_co_valid; // @[Core.scala 96:19:@24822.4]
  assign compute_io_inst_bits = fetch_io_inst_co_bits; // @[Core.scala 96:19:@24821.4]
  assign compute_io_uop_baddr = io_vcr_ptrs_1; // @[Core.scala 97:24:@24824.4]
  assign compute_io_acc_baddr = io_vcr_ptrs_4; // @[Core.scala 98:24:@24825.4]
  assign compute_io_vme_rd_0_cmd_ready = io_vme_rd_1_cmd_ready; // @[Core.scala 74:16:@24780.4]
  assign compute_io_vme_rd_0_data_valid = io_vme_rd_1_data_valid; // @[Core.scala 74:16:@24775.4]
  assign compute_io_vme_rd_0_data_bits = io_vme_rd_1_data_bits; // @[Core.scala 74:16:@24774.4]
  assign compute_io_vme_rd_1_cmd_ready = io_vme_rd_4_cmd_ready; // @[Core.scala 77:16:@24801.4]
  assign compute_io_vme_rd_1_data_valid = io_vme_rd_4_data_valid; // @[Core.scala 77:16:@24796.4]
  assign compute_io_vme_rd_1_data_bits = io_vme_rd_4_data_bits; // @[Core.scala 77:16:@24795.4]
  assign compute_io_inp_rd_data_valid = load_io_inp_rd_data_valid; // @[Core.scala 99:18:@24860.4]
  assign compute_io_inp_rd_data_bits_0_0 = load_io_inp_rd_data_bits_0_0; // @[Core.scala 99:18:@24844.4]
  assign compute_io_inp_rd_data_bits_0_1 = load_io_inp_rd_data_bits_0_1; // @[Core.scala 99:18:@24845.4]
  assign compute_io_inp_rd_data_bits_0_2 = load_io_inp_rd_data_bits_0_2; // @[Core.scala 99:18:@24846.4]
  assign compute_io_inp_rd_data_bits_0_3 = load_io_inp_rd_data_bits_0_3; // @[Core.scala 99:18:@24847.4]
  assign compute_io_inp_rd_data_bits_0_4 = load_io_inp_rd_data_bits_0_4; // @[Core.scala 99:18:@24848.4]
  assign compute_io_inp_rd_data_bits_0_5 = load_io_inp_rd_data_bits_0_5; // @[Core.scala 99:18:@24849.4]
  assign compute_io_inp_rd_data_bits_0_6 = load_io_inp_rd_data_bits_0_6; // @[Core.scala 99:18:@24850.4]
  assign compute_io_inp_rd_data_bits_0_7 = load_io_inp_rd_data_bits_0_7; // @[Core.scala 99:18:@24851.4]
  assign compute_io_inp_rd_data_bits_0_8 = load_io_inp_rd_data_bits_0_8; // @[Core.scala 99:18:@24852.4]
  assign compute_io_inp_rd_data_bits_0_9 = load_io_inp_rd_data_bits_0_9; // @[Core.scala 99:18:@24853.4]
  assign compute_io_inp_rd_data_bits_0_10 = load_io_inp_rd_data_bits_0_10; // @[Core.scala 99:18:@24854.4]
  assign compute_io_inp_rd_data_bits_0_11 = load_io_inp_rd_data_bits_0_11; // @[Core.scala 99:18:@24855.4]
  assign compute_io_inp_rd_data_bits_0_12 = load_io_inp_rd_data_bits_0_12; // @[Core.scala 99:18:@24856.4]
  assign compute_io_inp_rd_data_bits_0_13 = load_io_inp_rd_data_bits_0_13; // @[Core.scala 99:18:@24857.4]
  assign compute_io_inp_rd_data_bits_0_14 = load_io_inp_rd_data_bits_0_14; // @[Core.scala 99:18:@24858.4]
  assign compute_io_inp_rd_data_bits_0_15 = load_io_inp_rd_data_bits_0_15; // @[Core.scala 99:18:@24859.4]
  assign compute_io_wgt_rd_data_valid = load_io_wgt_rd_data_valid; // @[Core.scala 100:18:@25377.4]
  assign compute_io_wgt_rd_data_bits_0_0 = load_io_wgt_rd_data_bits_0_0; // @[Core.scala 100:18:@25121.4]
  assign compute_io_wgt_rd_data_bits_0_1 = load_io_wgt_rd_data_bits_0_1; // @[Core.scala 100:18:@25122.4]
  assign compute_io_wgt_rd_data_bits_0_2 = load_io_wgt_rd_data_bits_0_2; // @[Core.scala 100:18:@25123.4]
  assign compute_io_wgt_rd_data_bits_0_3 = load_io_wgt_rd_data_bits_0_3; // @[Core.scala 100:18:@25124.4]
  assign compute_io_wgt_rd_data_bits_0_4 = load_io_wgt_rd_data_bits_0_4; // @[Core.scala 100:18:@25125.4]
  assign compute_io_wgt_rd_data_bits_0_5 = load_io_wgt_rd_data_bits_0_5; // @[Core.scala 100:18:@25126.4]
  assign compute_io_wgt_rd_data_bits_0_6 = load_io_wgt_rd_data_bits_0_6; // @[Core.scala 100:18:@25127.4]
  assign compute_io_wgt_rd_data_bits_0_7 = load_io_wgt_rd_data_bits_0_7; // @[Core.scala 100:18:@25128.4]
  assign compute_io_wgt_rd_data_bits_0_8 = load_io_wgt_rd_data_bits_0_8; // @[Core.scala 100:18:@25129.4]
  assign compute_io_wgt_rd_data_bits_0_9 = load_io_wgt_rd_data_bits_0_9; // @[Core.scala 100:18:@25130.4]
  assign compute_io_wgt_rd_data_bits_0_10 = load_io_wgt_rd_data_bits_0_10; // @[Core.scala 100:18:@25131.4]
  assign compute_io_wgt_rd_data_bits_0_11 = load_io_wgt_rd_data_bits_0_11; // @[Core.scala 100:18:@25132.4]
  assign compute_io_wgt_rd_data_bits_0_12 = load_io_wgt_rd_data_bits_0_12; // @[Core.scala 100:18:@25133.4]
  assign compute_io_wgt_rd_data_bits_0_13 = load_io_wgt_rd_data_bits_0_13; // @[Core.scala 100:18:@25134.4]
  assign compute_io_wgt_rd_data_bits_0_14 = load_io_wgt_rd_data_bits_0_14; // @[Core.scala 100:18:@25135.4]
  assign compute_io_wgt_rd_data_bits_0_15 = load_io_wgt_rd_data_bits_0_15; // @[Core.scala 100:18:@25136.4]
  assign compute_io_wgt_rd_data_bits_1_0 = load_io_wgt_rd_data_bits_1_0; // @[Core.scala 100:18:@25137.4]
  assign compute_io_wgt_rd_data_bits_1_1 = load_io_wgt_rd_data_bits_1_1; // @[Core.scala 100:18:@25138.4]
  assign compute_io_wgt_rd_data_bits_1_2 = load_io_wgt_rd_data_bits_1_2; // @[Core.scala 100:18:@25139.4]
  assign compute_io_wgt_rd_data_bits_1_3 = load_io_wgt_rd_data_bits_1_3; // @[Core.scala 100:18:@25140.4]
  assign compute_io_wgt_rd_data_bits_1_4 = load_io_wgt_rd_data_bits_1_4; // @[Core.scala 100:18:@25141.4]
  assign compute_io_wgt_rd_data_bits_1_5 = load_io_wgt_rd_data_bits_1_5; // @[Core.scala 100:18:@25142.4]
  assign compute_io_wgt_rd_data_bits_1_6 = load_io_wgt_rd_data_bits_1_6; // @[Core.scala 100:18:@25143.4]
  assign compute_io_wgt_rd_data_bits_1_7 = load_io_wgt_rd_data_bits_1_7; // @[Core.scala 100:18:@25144.4]
  assign compute_io_wgt_rd_data_bits_1_8 = load_io_wgt_rd_data_bits_1_8; // @[Core.scala 100:18:@25145.4]
  assign compute_io_wgt_rd_data_bits_1_9 = load_io_wgt_rd_data_bits_1_9; // @[Core.scala 100:18:@25146.4]
  assign compute_io_wgt_rd_data_bits_1_10 = load_io_wgt_rd_data_bits_1_10; // @[Core.scala 100:18:@25147.4]
  assign compute_io_wgt_rd_data_bits_1_11 = load_io_wgt_rd_data_bits_1_11; // @[Core.scala 100:18:@25148.4]
  assign compute_io_wgt_rd_data_bits_1_12 = load_io_wgt_rd_data_bits_1_12; // @[Core.scala 100:18:@25149.4]
  assign compute_io_wgt_rd_data_bits_1_13 = load_io_wgt_rd_data_bits_1_13; // @[Core.scala 100:18:@25150.4]
  assign compute_io_wgt_rd_data_bits_1_14 = load_io_wgt_rd_data_bits_1_14; // @[Core.scala 100:18:@25151.4]
  assign compute_io_wgt_rd_data_bits_1_15 = load_io_wgt_rd_data_bits_1_15; // @[Core.scala 100:18:@25152.4]
  assign compute_io_wgt_rd_data_bits_2_0 = load_io_wgt_rd_data_bits_2_0; // @[Core.scala 100:18:@25153.4]
  assign compute_io_wgt_rd_data_bits_2_1 = load_io_wgt_rd_data_bits_2_1; // @[Core.scala 100:18:@25154.4]
  assign compute_io_wgt_rd_data_bits_2_2 = load_io_wgt_rd_data_bits_2_2; // @[Core.scala 100:18:@25155.4]
  assign compute_io_wgt_rd_data_bits_2_3 = load_io_wgt_rd_data_bits_2_3; // @[Core.scala 100:18:@25156.4]
  assign compute_io_wgt_rd_data_bits_2_4 = load_io_wgt_rd_data_bits_2_4; // @[Core.scala 100:18:@25157.4]
  assign compute_io_wgt_rd_data_bits_2_5 = load_io_wgt_rd_data_bits_2_5; // @[Core.scala 100:18:@25158.4]
  assign compute_io_wgt_rd_data_bits_2_6 = load_io_wgt_rd_data_bits_2_6; // @[Core.scala 100:18:@25159.4]
  assign compute_io_wgt_rd_data_bits_2_7 = load_io_wgt_rd_data_bits_2_7; // @[Core.scala 100:18:@25160.4]
  assign compute_io_wgt_rd_data_bits_2_8 = load_io_wgt_rd_data_bits_2_8; // @[Core.scala 100:18:@25161.4]
  assign compute_io_wgt_rd_data_bits_2_9 = load_io_wgt_rd_data_bits_2_9; // @[Core.scala 100:18:@25162.4]
  assign compute_io_wgt_rd_data_bits_2_10 = load_io_wgt_rd_data_bits_2_10; // @[Core.scala 100:18:@25163.4]
  assign compute_io_wgt_rd_data_bits_2_11 = load_io_wgt_rd_data_bits_2_11; // @[Core.scala 100:18:@25164.4]
  assign compute_io_wgt_rd_data_bits_2_12 = load_io_wgt_rd_data_bits_2_12; // @[Core.scala 100:18:@25165.4]
  assign compute_io_wgt_rd_data_bits_2_13 = load_io_wgt_rd_data_bits_2_13; // @[Core.scala 100:18:@25166.4]
  assign compute_io_wgt_rd_data_bits_2_14 = load_io_wgt_rd_data_bits_2_14; // @[Core.scala 100:18:@25167.4]
  assign compute_io_wgt_rd_data_bits_2_15 = load_io_wgt_rd_data_bits_2_15; // @[Core.scala 100:18:@25168.4]
  assign compute_io_wgt_rd_data_bits_3_0 = load_io_wgt_rd_data_bits_3_0; // @[Core.scala 100:18:@25169.4]
  assign compute_io_wgt_rd_data_bits_3_1 = load_io_wgt_rd_data_bits_3_1; // @[Core.scala 100:18:@25170.4]
  assign compute_io_wgt_rd_data_bits_3_2 = load_io_wgt_rd_data_bits_3_2; // @[Core.scala 100:18:@25171.4]
  assign compute_io_wgt_rd_data_bits_3_3 = load_io_wgt_rd_data_bits_3_3; // @[Core.scala 100:18:@25172.4]
  assign compute_io_wgt_rd_data_bits_3_4 = load_io_wgt_rd_data_bits_3_4; // @[Core.scala 100:18:@25173.4]
  assign compute_io_wgt_rd_data_bits_3_5 = load_io_wgt_rd_data_bits_3_5; // @[Core.scala 100:18:@25174.4]
  assign compute_io_wgt_rd_data_bits_3_6 = load_io_wgt_rd_data_bits_3_6; // @[Core.scala 100:18:@25175.4]
  assign compute_io_wgt_rd_data_bits_3_7 = load_io_wgt_rd_data_bits_3_7; // @[Core.scala 100:18:@25176.4]
  assign compute_io_wgt_rd_data_bits_3_8 = load_io_wgt_rd_data_bits_3_8; // @[Core.scala 100:18:@25177.4]
  assign compute_io_wgt_rd_data_bits_3_9 = load_io_wgt_rd_data_bits_3_9; // @[Core.scala 100:18:@25178.4]
  assign compute_io_wgt_rd_data_bits_3_10 = load_io_wgt_rd_data_bits_3_10; // @[Core.scala 100:18:@25179.4]
  assign compute_io_wgt_rd_data_bits_3_11 = load_io_wgt_rd_data_bits_3_11; // @[Core.scala 100:18:@25180.4]
  assign compute_io_wgt_rd_data_bits_3_12 = load_io_wgt_rd_data_bits_3_12; // @[Core.scala 100:18:@25181.4]
  assign compute_io_wgt_rd_data_bits_3_13 = load_io_wgt_rd_data_bits_3_13; // @[Core.scala 100:18:@25182.4]
  assign compute_io_wgt_rd_data_bits_3_14 = load_io_wgt_rd_data_bits_3_14; // @[Core.scala 100:18:@25183.4]
  assign compute_io_wgt_rd_data_bits_3_15 = load_io_wgt_rd_data_bits_3_15; // @[Core.scala 100:18:@25184.4]
  assign compute_io_wgt_rd_data_bits_4_0 = load_io_wgt_rd_data_bits_4_0; // @[Core.scala 100:18:@25185.4]
  assign compute_io_wgt_rd_data_bits_4_1 = load_io_wgt_rd_data_bits_4_1; // @[Core.scala 100:18:@25186.4]
  assign compute_io_wgt_rd_data_bits_4_2 = load_io_wgt_rd_data_bits_4_2; // @[Core.scala 100:18:@25187.4]
  assign compute_io_wgt_rd_data_bits_4_3 = load_io_wgt_rd_data_bits_4_3; // @[Core.scala 100:18:@25188.4]
  assign compute_io_wgt_rd_data_bits_4_4 = load_io_wgt_rd_data_bits_4_4; // @[Core.scala 100:18:@25189.4]
  assign compute_io_wgt_rd_data_bits_4_5 = load_io_wgt_rd_data_bits_4_5; // @[Core.scala 100:18:@25190.4]
  assign compute_io_wgt_rd_data_bits_4_6 = load_io_wgt_rd_data_bits_4_6; // @[Core.scala 100:18:@25191.4]
  assign compute_io_wgt_rd_data_bits_4_7 = load_io_wgt_rd_data_bits_4_7; // @[Core.scala 100:18:@25192.4]
  assign compute_io_wgt_rd_data_bits_4_8 = load_io_wgt_rd_data_bits_4_8; // @[Core.scala 100:18:@25193.4]
  assign compute_io_wgt_rd_data_bits_4_9 = load_io_wgt_rd_data_bits_4_9; // @[Core.scala 100:18:@25194.4]
  assign compute_io_wgt_rd_data_bits_4_10 = load_io_wgt_rd_data_bits_4_10; // @[Core.scala 100:18:@25195.4]
  assign compute_io_wgt_rd_data_bits_4_11 = load_io_wgt_rd_data_bits_4_11; // @[Core.scala 100:18:@25196.4]
  assign compute_io_wgt_rd_data_bits_4_12 = load_io_wgt_rd_data_bits_4_12; // @[Core.scala 100:18:@25197.4]
  assign compute_io_wgt_rd_data_bits_4_13 = load_io_wgt_rd_data_bits_4_13; // @[Core.scala 100:18:@25198.4]
  assign compute_io_wgt_rd_data_bits_4_14 = load_io_wgt_rd_data_bits_4_14; // @[Core.scala 100:18:@25199.4]
  assign compute_io_wgt_rd_data_bits_4_15 = load_io_wgt_rd_data_bits_4_15; // @[Core.scala 100:18:@25200.4]
  assign compute_io_wgt_rd_data_bits_5_0 = load_io_wgt_rd_data_bits_5_0; // @[Core.scala 100:18:@25201.4]
  assign compute_io_wgt_rd_data_bits_5_1 = load_io_wgt_rd_data_bits_5_1; // @[Core.scala 100:18:@25202.4]
  assign compute_io_wgt_rd_data_bits_5_2 = load_io_wgt_rd_data_bits_5_2; // @[Core.scala 100:18:@25203.4]
  assign compute_io_wgt_rd_data_bits_5_3 = load_io_wgt_rd_data_bits_5_3; // @[Core.scala 100:18:@25204.4]
  assign compute_io_wgt_rd_data_bits_5_4 = load_io_wgt_rd_data_bits_5_4; // @[Core.scala 100:18:@25205.4]
  assign compute_io_wgt_rd_data_bits_5_5 = load_io_wgt_rd_data_bits_5_5; // @[Core.scala 100:18:@25206.4]
  assign compute_io_wgt_rd_data_bits_5_6 = load_io_wgt_rd_data_bits_5_6; // @[Core.scala 100:18:@25207.4]
  assign compute_io_wgt_rd_data_bits_5_7 = load_io_wgt_rd_data_bits_5_7; // @[Core.scala 100:18:@25208.4]
  assign compute_io_wgt_rd_data_bits_5_8 = load_io_wgt_rd_data_bits_5_8; // @[Core.scala 100:18:@25209.4]
  assign compute_io_wgt_rd_data_bits_5_9 = load_io_wgt_rd_data_bits_5_9; // @[Core.scala 100:18:@25210.4]
  assign compute_io_wgt_rd_data_bits_5_10 = load_io_wgt_rd_data_bits_5_10; // @[Core.scala 100:18:@25211.4]
  assign compute_io_wgt_rd_data_bits_5_11 = load_io_wgt_rd_data_bits_5_11; // @[Core.scala 100:18:@25212.4]
  assign compute_io_wgt_rd_data_bits_5_12 = load_io_wgt_rd_data_bits_5_12; // @[Core.scala 100:18:@25213.4]
  assign compute_io_wgt_rd_data_bits_5_13 = load_io_wgt_rd_data_bits_5_13; // @[Core.scala 100:18:@25214.4]
  assign compute_io_wgt_rd_data_bits_5_14 = load_io_wgt_rd_data_bits_5_14; // @[Core.scala 100:18:@25215.4]
  assign compute_io_wgt_rd_data_bits_5_15 = load_io_wgt_rd_data_bits_5_15; // @[Core.scala 100:18:@25216.4]
  assign compute_io_wgt_rd_data_bits_6_0 = load_io_wgt_rd_data_bits_6_0; // @[Core.scala 100:18:@25217.4]
  assign compute_io_wgt_rd_data_bits_6_1 = load_io_wgt_rd_data_bits_6_1; // @[Core.scala 100:18:@25218.4]
  assign compute_io_wgt_rd_data_bits_6_2 = load_io_wgt_rd_data_bits_6_2; // @[Core.scala 100:18:@25219.4]
  assign compute_io_wgt_rd_data_bits_6_3 = load_io_wgt_rd_data_bits_6_3; // @[Core.scala 100:18:@25220.4]
  assign compute_io_wgt_rd_data_bits_6_4 = load_io_wgt_rd_data_bits_6_4; // @[Core.scala 100:18:@25221.4]
  assign compute_io_wgt_rd_data_bits_6_5 = load_io_wgt_rd_data_bits_6_5; // @[Core.scala 100:18:@25222.4]
  assign compute_io_wgt_rd_data_bits_6_6 = load_io_wgt_rd_data_bits_6_6; // @[Core.scala 100:18:@25223.4]
  assign compute_io_wgt_rd_data_bits_6_7 = load_io_wgt_rd_data_bits_6_7; // @[Core.scala 100:18:@25224.4]
  assign compute_io_wgt_rd_data_bits_6_8 = load_io_wgt_rd_data_bits_6_8; // @[Core.scala 100:18:@25225.4]
  assign compute_io_wgt_rd_data_bits_6_9 = load_io_wgt_rd_data_bits_6_9; // @[Core.scala 100:18:@25226.4]
  assign compute_io_wgt_rd_data_bits_6_10 = load_io_wgt_rd_data_bits_6_10; // @[Core.scala 100:18:@25227.4]
  assign compute_io_wgt_rd_data_bits_6_11 = load_io_wgt_rd_data_bits_6_11; // @[Core.scala 100:18:@25228.4]
  assign compute_io_wgt_rd_data_bits_6_12 = load_io_wgt_rd_data_bits_6_12; // @[Core.scala 100:18:@25229.4]
  assign compute_io_wgt_rd_data_bits_6_13 = load_io_wgt_rd_data_bits_6_13; // @[Core.scala 100:18:@25230.4]
  assign compute_io_wgt_rd_data_bits_6_14 = load_io_wgt_rd_data_bits_6_14; // @[Core.scala 100:18:@25231.4]
  assign compute_io_wgt_rd_data_bits_6_15 = load_io_wgt_rd_data_bits_6_15; // @[Core.scala 100:18:@25232.4]
  assign compute_io_wgt_rd_data_bits_7_0 = load_io_wgt_rd_data_bits_7_0; // @[Core.scala 100:18:@25233.4]
  assign compute_io_wgt_rd_data_bits_7_1 = load_io_wgt_rd_data_bits_7_1; // @[Core.scala 100:18:@25234.4]
  assign compute_io_wgt_rd_data_bits_7_2 = load_io_wgt_rd_data_bits_7_2; // @[Core.scala 100:18:@25235.4]
  assign compute_io_wgt_rd_data_bits_7_3 = load_io_wgt_rd_data_bits_7_3; // @[Core.scala 100:18:@25236.4]
  assign compute_io_wgt_rd_data_bits_7_4 = load_io_wgt_rd_data_bits_7_4; // @[Core.scala 100:18:@25237.4]
  assign compute_io_wgt_rd_data_bits_7_5 = load_io_wgt_rd_data_bits_7_5; // @[Core.scala 100:18:@25238.4]
  assign compute_io_wgt_rd_data_bits_7_6 = load_io_wgt_rd_data_bits_7_6; // @[Core.scala 100:18:@25239.4]
  assign compute_io_wgt_rd_data_bits_7_7 = load_io_wgt_rd_data_bits_7_7; // @[Core.scala 100:18:@25240.4]
  assign compute_io_wgt_rd_data_bits_7_8 = load_io_wgt_rd_data_bits_7_8; // @[Core.scala 100:18:@25241.4]
  assign compute_io_wgt_rd_data_bits_7_9 = load_io_wgt_rd_data_bits_7_9; // @[Core.scala 100:18:@25242.4]
  assign compute_io_wgt_rd_data_bits_7_10 = load_io_wgt_rd_data_bits_7_10; // @[Core.scala 100:18:@25243.4]
  assign compute_io_wgt_rd_data_bits_7_11 = load_io_wgt_rd_data_bits_7_11; // @[Core.scala 100:18:@25244.4]
  assign compute_io_wgt_rd_data_bits_7_12 = load_io_wgt_rd_data_bits_7_12; // @[Core.scala 100:18:@25245.4]
  assign compute_io_wgt_rd_data_bits_7_13 = load_io_wgt_rd_data_bits_7_13; // @[Core.scala 100:18:@25246.4]
  assign compute_io_wgt_rd_data_bits_7_14 = load_io_wgt_rd_data_bits_7_14; // @[Core.scala 100:18:@25247.4]
  assign compute_io_wgt_rd_data_bits_7_15 = load_io_wgt_rd_data_bits_7_15; // @[Core.scala 100:18:@25248.4]
  assign compute_io_wgt_rd_data_bits_8_0 = load_io_wgt_rd_data_bits_8_0; // @[Core.scala 100:18:@25249.4]
  assign compute_io_wgt_rd_data_bits_8_1 = load_io_wgt_rd_data_bits_8_1; // @[Core.scala 100:18:@25250.4]
  assign compute_io_wgt_rd_data_bits_8_2 = load_io_wgt_rd_data_bits_8_2; // @[Core.scala 100:18:@25251.4]
  assign compute_io_wgt_rd_data_bits_8_3 = load_io_wgt_rd_data_bits_8_3; // @[Core.scala 100:18:@25252.4]
  assign compute_io_wgt_rd_data_bits_8_4 = load_io_wgt_rd_data_bits_8_4; // @[Core.scala 100:18:@25253.4]
  assign compute_io_wgt_rd_data_bits_8_5 = load_io_wgt_rd_data_bits_8_5; // @[Core.scala 100:18:@25254.4]
  assign compute_io_wgt_rd_data_bits_8_6 = load_io_wgt_rd_data_bits_8_6; // @[Core.scala 100:18:@25255.4]
  assign compute_io_wgt_rd_data_bits_8_7 = load_io_wgt_rd_data_bits_8_7; // @[Core.scala 100:18:@25256.4]
  assign compute_io_wgt_rd_data_bits_8_8 = load_io_wgt_rd_data_bits_8_8; // @[Core.scala 100:18:@25257.4]
  assign compute_io_wgt_rd_data_bits_8_9 = load_io_wgt_rd_data_bits_8_9; // @[Core.scala 100:18:@25258.4]
  assign compute_io_wgt_rd_data_bits_8_10 = load_io_wgt_rd_data_bits_8_10; // @[Core.scala 100:18:@25259.4]
  assign compute_io_wgt_rd_data_bits_8_11 = load_io_wgt_rd_data_bits_8_11; // @[Core.scala 100:18:@25260.4]
  assign compute_io_wgt_rd_data_bits_8_12 = load_io_wgt_rd_data_bits_8_12; // @[Core.scala 100:18:@25261.4]
  assign compute_io_wgt_rd_data_bits_8_13 = load_io_wgt_rd_data_bits_8_13; // @[Core.scala 100:18:@25262.4]
  assign compute_io_wgt_rd_data_bits_8_14 = load_io_wgt_rd_data_bits_8_14; // @[Core.scala 100:18:@25263.4]
  assign compute_io_wgt_rd_data_bits_8_15 = load_io_wgt_rd_data_bits_8_15; // @[Core.scala 100:18:@25264.4]
  assign compute_io_wgt_rd_data_bits_9_0 = load_io_wgt_rd_data_bits_9_0; // @[Core.scala 100:18:@25265.4]
  assign compute_io_wgt_rd_data_bits_9_1 = load_io_wgt_rd_data_bits_9_1; // @[Core.scala 100:18:@25266.4]
  assign compute_io_wgt_rd_data_bits_9_2 = load_io_wgt_rd_data_bits_9_2; // @[Core.scala 100:18:@25267.4]
  assign compute_io_wgt_rd_data_bits_9_3 = load_io_wgt_rd_data_bits_9_3; // @[Core.scala 100:18:@25268.4]
  assign compute_io_wgt_rd_data_bits_9_4 = load_io_wgt_rd_data_bits_9_4; // @[Core.scala 100:18:@25269.4]
  assign compute_io_wgt_rd_data_bits_9_5 = load_io_wgt_rd_data_bits_9_5; // @[Core.scala 100:18:@25270.4]
  assign compute_io_wgt_rd_data_bits_9_6 = load_io_wgt_rd_data_bits_9_6; // @[Core.scala 100:18:@25271.4]
  assign compute_io_wgt_rd_data_bits_9_7 = load_io_wgt_rd_data_bits_9_7; // @[Core.scala 100:18:@25272.4]
  assign compute_io_wgt_rd_data_bits_9_8 = load_io_wgt_rd_data_bits_9_8; // @[Core.scala 100:18:@25273.4]
  assign compute_io_wgt_rd_data_bits_9_9 = load_io_wgt_rd_data_bits_9_9; // @[Core.scala 100:18:@25274.4]
  assign compute_io_wgt_rd_data_bits_9_10 = load_io_wgt_rd_data_bits_9_10; // @[Core.scala 100:18:@25275.4]
  assign compute_io_wgt_rd_data_bits_9_11 = load_io_wgt_rd_data_bits_9_11; // @[Core.scala 100:18:@25276.4]
  assign compute_io_wgt_rd_data_bits_9_12 = load_io_wgt_rd_data_bits_9_12; // @[Core.scala 100:18:@25277.4]
  assign compute_io_wgt_rd_data_bits_9_13 = load_io_wgt_rd_data_bits_9_13; // @[Core.scala 100:18:@25278.4]
  assign compute_io_wgt_rd_data_bits_9_14 = load_io_wgt_rd_data_bits_9_14; // @[Core.scala 100:18:@25279.4]
  assign compute_io_wgt_rd_data_bits_9_15 = load_io_wgt_rd_data_bits_9_15; // @[Core.scala 100:18:@25280.4]
  assign compute_io_wgt_rd_data_bits_10_0 = load_io_wgt_rd_data_bits_10_0; // @[Core.scala 100:18:@25281.4]
  assign compute_io_wgt_rd_data_bits_10_1 = load_io_wgt_rd_data_bits_10_1; // @[Core.scala 100:18:@25282.4]
  assign compute_io_wgt_rd_data_bits_10_2 = load_io_wgt_rd_data_bits_10_2; // @[Core.scala 100:18:@25283.4]
  assign compute_io_wgt_rd_data_bits_10_3 = load_io_wgt_rd_data_bits_10_3; // @[Core.scala 100:18:@25284.4]
  assign compute_io_wgt_rd_data_bits_10_4 = load_io_wgt_rd_data_bits_10_4; // @[Core.scala 100:18:@25285.4]
  assign compute_io_wgt_rd_data_bits_10_5 = load_io_wgt_rd_data_bits_10_5; // @[Core.scala 100:18:@25286.4]
  assign compute_io_wgt_rd_data_bits_10_6 = load_io_wgt_rd_data_bits_10_6; // @[Core.scala 100:18:@25287.4]
  assign compute_io_wgt_rd_data_bits_10_7 = load_io_wgt_rd_data_bits_10_7; // @[Core.scala 100:18:@25288.4]
  assign compute_io_wgt_rd_data_bits_10_8 = load_io_wgt_rd_data_bits_10_8; // @[Core.scala 100:18:@25289.4]
  assign compute_io_wgt_rd_data_bits_10_9 = load_io_wgt_rd_data_bits_10_9; // @[Core.scala 100:18:@25290.4]
  assign compute_io_wgt_rd_data_bits_10_10 = load_io_wgt_rd_data_bits_10_10; // @[Core.scala 100:18:@25291.4]
  assign compute_io_wgt_rd_data_bits_10_11 = load_io_wgt_rd_data_bits_10_11; // @[Core.scala 100:18:@25292.4]
  assign compute_io_wgt_rd_data_bits_10_12 = load_io_wgt_rd_data_bits_10_12; // @[Core.scala 100:18:@25293.4]
  assign compute_io_wgt_rd_data_bits_10_13 = load_io_wgt_rd_data_bits_10_13; // @[Core.scala 100:18:@25294.4]
  assign compute_io_wgt_rd_data_bits_10_14 = load_io_wgt_rd_data_bits_10_14; // @[Core.scala 100:18:@25295.4]
  assign compute_io_wgt_rd_data_bits_10_15 = load_io_wgt_rd_data_bits_10_15; // @[Core.scala 100:18:@25296.4]
  assign compute_io_wgt_rd_data_bits_11_0 = load_io_wgt_rd_data_bits_11_0; // @[Core.scala 100:18:@25297.4]
  assign compute_io_wgt_rd_data_bits_11_1 = load_io_wgt_rd_data_bits_11_1; // @[Core.scala 100:18:@25298.4]
  assign compute_io_wgt_rd_data_bits_11_2 = load_io_wgt_rd_data_bits_11_2; // @[Core.scala 100:18:@25299.4]
  assign compute_io_wgt_rd_data_bits_11_3 = load_io_wgt_rd_data_bits_11_3; // @[Core.scala 100:18:@25300.4]
  assign compute_io_wgt_rd_data_bits_11_4 = load_io_wgt_rd_data_bits_11_4; // @[Core.scala 100:18:@25301.4]
  assign compute_io_wgt_rd_data_bits_11_5 = load_io_wgt_rd_data_bits_11_5; // @[Core.scala 100:18:@25302.4]
  assign compute_io_wgt_rd_data_bits_11_6 = load_io_wgt_rd_data_bits_11_6; // @[Core.scala 100:18:@25303.4]
  assign compute_io_wgt_rd_data_bits_11_7 = load_io_wgt_rd_data_bits_11_7; // @[Core.scala 100:18:@25304.4]
  assign compute_io_wgt_rd_data_bits_11_8 = load_io_wgt_rd_data_bits_11_8; // @[Core.scala 100:18:@25305.4]
  assign compute_io_wgt_rd_data_bits_11_9 = load_io_wgt_rd_data_bits_11_9; // @[Core.scala 100:18:@25306.4]
  assign compute_io_wgt_rd_data_bits_11_10 = load_io_wgt_rd_data_bits_11_10; // @[Core.scala 100:18:@25307.4]
  assign compute_io_wgt_rd_data_bits_11_11 = load_io_wgt_rd_data_bits_11_11; // @[Core.scala 100:18:@25308.4]
  assign compute_io_wgt_rd_data_bits_11_12 = load_io_wgt_rd_data_bits_11_12; // @[Core.scala 100:18:@25309.4]
  assign compute_io_wgt_rd_data_bits_11_13 = load_io_wgt_rd_data_bits_11_13; // @[Core.scala 100:18:@25310.4]
  assign compute_io_wgt_rd_data_bits_11_14 = load_io_wgt_rd_data_bits_11_14; // @[Core.scala 100:18:@25311.4]
  assign compute_io_wgt_rd_data_bits_11_15 = load_io_wgt_rd_data_bits_11_15; // @[Core.scala 100:18:@25312.4]
  assign compute_io_wgt_rd_data_bits_12_0 = load_io_wgt_rd_data_bits_12_0; // @[Core.scala 100:18:@25313.4]
  assign compute_io_wgt_rd_data_bits_12_1 = load_io_wgt_rd_data_bits_12_1; // @[Core.scala 100:18:@25314.4]
  assign compute_io_wgt_rd_data_bits_12_2 = load_io_wgt_rd_data_bits_12_2; // @[Core.scala 100:18:@25315.4]
  assign compute_io_wgt_rd_data_bits_12_3 = load_io_wgt_rd_data_bits_12_3; // @[Core.scala 100:18:@25316.4]
  assign compute_io_wgt_rd_data_bits_12_4 = load_io_wgt_rd_data_bits_12_4; // @[Core.scala 100:18:@25317.4]
  assign compute_io_wgt_rd_data_bits_12_5 = load_io_wgt_rd_data_bits_12_5; // @[Core.scala 100:18:@25318.4]
  assign compute_io_wgt_rd_data_bits_12_6 = load_io_wgt_rd_data_bits_12_6; // @[Core.scala 100:18:@25319.4]
  assign compute_io_wgt_rd_data_bits_12_7 = load_io_wgt_rd_data_bits_12_7; // @[Core.scala 100:18:@25320.4]
  assign compute_io_wgt_rd_data_bits_12_8 = load_io_wgt_rd_data_bits_12_8; // @[Core.scala 100:18:@25321.4]
  assign compute_io_wgt_rd_data_bits_12_9 = load_io_wgt_rd_data_bits_12_9; // @[Core.scala 100:18:@25322.4]
  assign compute_io_wgt_rd_data_bits_12_10 = load_io_wgt_rd_data_bits_12_10; // @[Core.scala 100:18:@25323.4]
  assign compute_io_wgt_rd_data_bits_12_11 = load_io_wgt_rd_data_bits_12_11; // @[Core.scala 100:18:@25324.4]
  assign compute_io_wgt_rd_data_bits_12_12 = load_io_wgt_rd_data_bits_12_12; // @[Core.scala 100:18:@25325.4]
  assign compute_io_wgt_rd_data_bits_12_13 = load_io_wgt_rd_data_bits_12_13; // @[Core.scala 100:18:@25326.4]
  assign compute_io_wgt_rd_data_bits_12_14 = load_io_wgt_rd_data_bits_12_14; // @[Core.scala 100:18:@25327.4]
  assign compute_io_wgt_rd_data_bits_12_15 = load_io_wgt_rd_data_bits_12_15; // @[Core.scala 100:18:@25328.4]
  assign compute_io_wgt_rd_data_bits_13_0 = load_io_wgt_rd_data_bits_13_0; // @[Core.scala 100:18:@25329.4]
  assign compute_io_wgt_rd_data_bits_13_1 = load_io_wgt_rd_data_bits_13_1; // @[Core.scala 100:18:@25330.4]
  assign compute_io_wgt_rd_data_bits_13_2 = load_io_wgt_rd_data_bits_13_2; // @[Core.scala 100:18:@25331.4]
  assign compute_io_wgt_rd_data_bits_13_3 = load_io_wgt_rd_data_bits_13_3; // @[Core.scala 100:18:@25332.4]
  assign compute_io_wgt_rd_data_bits_13_4 = load_io_wgt_rd_data_bits_13_4; // @[Core.scala 100:18:@25333.4]
  assign compute_io_wgt_rd_data_bits_13_5 = load_io_wgt_rd_data_bits_13_5; // @[Core.scala 100:18:@25334.4]
  assign compute_io_wgt_rd_data_bits_13_6 = load_io_wgt_rd_data_bits_13_6; // @[Core.scala 100:18:@25335.4]
  assign compute_io_wgt_rd_data_bits_13_7 = load_io_wgt_rd_data_bits_13_7; // @[Core.scala 100:18:@25336.4]
  assign compute_io_wgt_rd_data_bits_13_8 = load_io_wgt_rd_data_bits_13_8; // @[Core.scala 100:18:@25337.4]
  assign compute_io_wgt_rd_data_bits_13_9 = load_io_wgt_rd_data_bits_13_9; // @[Core.scala 100:18:@25338.4]
  assign compute_io_wgt_rd_data_bits_13_10 = load_io_wgt_rd_data_bits_13_10; // @[Core.scala 100:18:@25339.4]
  assign compute_io_wgt_rd_data_bits_13_11 = load_io_wgt_rd_data_bits_13_11; // @[Core.scala 100:18:@25340.4]
  assign compute_io_wgt_rd_data_bits_13_12 = load_io_wgt_rd_data_bits_13_12; // @[Core.scala 100:18:@25341.4]
  assign compute_io_wgt_rd_data_bits_13_13 = load_io_wgt_rd_data_bits_13_13; // @[Core.scala 100:18:@25342.4]
  assign compute_io_wgt_rd_data_bits_13_14 = load_io_wgt_rd_data_bits_13_14; // @[Core.scala 100:18:@25343.4]
  assign compute_io_wgt_rd_data_bits_13_15 = load_io_wgt_rd_data_bits_13_15; // @[Core.scala 100:18:@25344.4]
  assign compute_io_wgt_rd_data_bits_14_0 = load_io_wgt_rd_data_bits_14_0; // @[Core.scala 100:18:@25345.4]
  assign compute_io_wgt_rd_data_bits_14_1 = load_io_wgt_rd_data_bits_14_1; // @[Core.scala 100:18:@25346.4]
  assign compute_io_wgt_rd_data_bits_14_2 = load_io_wgt_rd_data_bits_14_2; // @[Core.scala 100:18:@25347.4]
  assign compute_io_wgt_rd_data_bits_14_3 = load_io_wgt_rd_data_bits_14_3; // @[Core.scala 100:18:@25348.4]
  assign compute_io_wgt_rd_data_bits_14_4 = load_io_wgt_rd_data_bits_14_4; // @[Core.scala 100:18:@25349.4]
  assign compute_io_wgt_rd_data_bits_14_5 = load_io_wgt_rd_data_bits_14_5; // @[Core.scala 100:18:@25350.4]
  assign compute_io_wgt_rd_data_bits_14_6 = load_io_wgt_rd_data_bits_14_6; // @[Core.scala 100:18:@25351.4]
  assign compute_io_wgt_rd_data_bits_14_7 = load_io_wgt_rd_data_bits_14_7; // @[Core.scala 100:18:@25352.4]
  assign compute_io_wgt_rd_data_bits_14_8 = load_io_wgt_rd_data_bits_14_8; // @[Core.scala 100:18:@25353.4]
  assign compute_io_wgt_rd_data_bits_14_9 = load_io_wgt_rd_data_bits_14_9; // @[Core.scala 100:18:@25354.4]
  assign compute_io_wgt_rd_data_bits_14_10 = load_io_wgt_rd_data_bits_14_10; // @[Core.scala 100:18:@25355.4]
  assign compute_io_wgt_rd_data_bits_14_11 = load_io_wgt_rd_data_bits_14_11; // @[Core.scala 100:18:@25356.4]
  assign compute_io_wgt_rd_data_bits_14_12 = load_io_wgt_rd_data_bits_14_12; // @[Core.scala 100:18:@25357.4]
  assign compute_io_wgt_rd_data_bits_14_13 = load_io_wgt_rd_data_bits_14_13; // @[Core.scala 100:18:@25358.4]
  assign compute_io_wgt_rd_data_bits_14_14 = load_io_wgt_rd_data_bits_14_14; // @[Core.scala 100:18:@25359.4]
  assign compute_io_wgt_rd_data_bits_14_15 = load_io_wgt_rd_data_bits_14_15; // @[Core.scala 100:18:@25360.4]
  assign compute_io_wgt_rd_data_bits_15_0 = load_io_wgt_rd_data_bits_15_0; // @[Core.scala 100:18:@25361.4]
  assign compute_io_wgt_rd_data_bits_15_1 = load_io_wgt_rd_data_bits_15_1; // @[Core.scala 100:18:@25362.4]
  assign compute_io_wgt_rd_data_bits_15_2 = load_io_wgt_rd_data_bits_15_2; // @[Core.scala 100:18:@25363.4]
  assign compute_io_wgt_rd_data_bits_15_3 = load_io_wgt_rd_data_bits_15_3; // @[Core.scala 100:18:@25364.4]
  assign compute_io_wgt_rd_data_bits_15_4 = load_io_wgt_rd_data_bits_15_4; // @[Core.scala 100:18:@25365.4]
  assign compute_io_wgt_rd_data_bits_15_5 = load_io_wgt_rd_data_bits_15_5; // @[Core.scala 100:18:@25366.4]
  assign compute_io_wgt_rd_data_bits_15_6 = load_io_wgt_rd_data_bits_15_6; // @[Core.scala 100:18:@25367.4]
  assign compute_io_wgt_rd_data_bits_15_7 = load_io_wgt_rd_data_bits_15_7; // @[Core.scala 100:18:@25368.4]
  assign compute_io_wgt_rd_data_bits_15_8 = load_io_wgt_rd_data_bits_15_8; // @[Core.scala 100:18:@25369.4]
  assign compute_io_wgt_rd_data_bits_15_9 = load_io_wgt_rd_data_bits_15_9; // @[Core.scala 100:18:@25370.4]
  assign compute_io_wgt_rd_data_bits_15_10 = load_io_wgt_rd_data_bits_15_10; // @[Core.scala 100:18:@25371.4]
  assign compute_io_wgt_rd_data_bits_15_11 = load_io_wgt_rd_data_bits_15_11; // @[Core.scala 100:18:@25372.4]
  assign compute_io_wgt_rd_data_bits_15_12 = load_io_wgt_rd_data_bits_15_12; // @[Core.scala 100:18:@25373.4]
  assign compute_io_wgt_rd_data_bits_15_13 = load_io_wgt_rd_data_bits_15_13; // @[Core.scala 100:18:@25374.4]
  assign compute_io_wgt_rd_data_bits_15_14 = load_io_wgt_rd_data_bits_15_14; // @[Core.scala 100:18:@25375.4]
  assign compute_io_wgt_rd_data_bits_15_15 = load_io_wgt_rd_data_bits_15_15; // @[Core.scala 100:18:@25376.4]
  assign store_clock = clock; // @[:@24762.4]
  assign store_reset = reset; // @[:@24763.4]
  assign store_io_i_post = compute_io_o_post_1; // @[Core.scala 105:19:@25380.4]
  assign store_io_inst_valid = fetch_io_inst_st_valid; // @[Core.scala 106:17:@25382.4]
  assign store_io_inst_bits = fetch_io_inst_st_bits; // @[Core.scala 106:17:@25381.4]
  assign store_io_out_baddr = io_vcr_ptrs_5; // @[Core.scala 107:22:@25384.4]
  assign store_io_vme_wr_cmd_ready = io_vme_wr_0_cmd_ready; // @[Core.scala 78:16:@24809.4]
  assign store_io_vme_wr_data_ready = io_vme_wr_0_data_ready; // @[Core.scala 78:16:@24805.4]
  assign store_io_vme_wr_ack = io_vme_wr_0_ack; // @[Core.scala 78:16:@24802.4]
  assign store_io_out_wr_valid = compute_io_out_wr_valid; // @[Core.scala 108:16:@25402.4]
  assign store_io_out_wr_bits_idx = compute_io_out_wr_bits_idx; // @[Core.scala 108:16:@25401.4]
  assign store_io_out_wr_bits_data_0_0 = compute_io_out_wr_bits_data_0_0; // @[Core.scala 108:16:@25385.4]
  assign store_io_out_wr_bits_data_0_1 = compute_io_out_wr_bits_data_0_1; // @[Core.scala 108:16:@25386.4]
  assign store_io_out_wr_bits_data_0_2 = compute_io_out_wr_bits_data_0_2; // @[Core.scala 108:16:@25387.4]
  assign store_io_out_wr_bits_data_0_3 = compute_io_out_wr_bits_data_0_3; // @[Core.scala 108:16:@25388.4]
  assign store_io_out_wr_bits_data_0_4 = compute_io_out_wr_bits_data_0_4; // @[Core.scala 108:16:@25389.4]
  assign store_io_out_wr_bits_data_0_5 = compute_io_out_wr_bits_data_0_5; // @[Core.scala 108:16:@25390.4]
  assign store_io_out_wr_bits_data_0_6 = compute_io_out_wr_bits_data_0_6; // @[Core.scala 108:16:@25391.4]
  assign store_io_out_wr_bits_data_0_7 = compute_io_out_wr_bits_data_0_7; // @[Core.scala 108:16:@25392.4]
  assign store_io_out_wr_bits_data_0_8 = compute_io_out_wr_bits_data_0_8; // @[Core.scala 108:16:@25393.4]
  assign store_io_out_wr_bits_data_0_9 = compute_io_out_wr_bits_data_0_9; // @[Core.scala 108:16:@25394.4]
  assign store_io_out_wr_bits_data_0_10 = compute_io_out_wr_bits_data_0_10; // @[Core.scala 108:16:@25395.4]
  assign store_io_out_wr_bits_data_0_11 = compute_io_out_wr_bits_data_0_11; // @[Core.scala 108:16:@25396.4]
  assign store_io_out_wr_bits_data_0_12 = compute_io_out_wr_bits_data_0_12; // @[Core.scala 108:16:@25397.4]
  assign store_io_out_wr_bits_data_0_13 = compute_io_out_wr_bits_data_0_13; // @[Core.scala 108:16:@25398.4]
  assign store_io_out_wr_bits_data_0_14 = compute_io_out_wr_bits_data_0_14; // @[Core.scala 108:16:@25399.4]
  assign store_io_out_wr_bits_data_0_15 = compute_io_out_wr_bits_data_0_15; // @[Core.scala 108:16:@25400.4]
  assign ecounters_clock = clock; // @[:@24765.4]
  assign ecounters_reset = reset; // @[:@24766.4]
  assign ecounters_io_launch = io_vcr_launch; // @[Core.scala 111:23:@25422.4]
  assign ecounters_io_finish = compute_io_finish; // @[Core.scala 112:23:@25423.4]
  assign ecounters_io_acc_wr_event = compute_io_acc_wr_event; // @[Core.scala 115:29:@25428.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  finish = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    finish <= compute_io_finish;
  end
endmodule
module VTAShell( // @[:@25433.2]
  input         clock, // @[:@25434.4]
  input         reset, // @[:@25435.4]
  output        io_host_aw_ready, // @[:@25436.4]
  input         io_host_aw_valid, // @[:@25436.4]
  input  [15:0] io_host_aw_bits_addr, // @[:@25436.4]
  output        io_host_w_ready, // @[:@25436.4]
  input         io_host_w_valid, // @[:@25436.4]
  input  [31:0] io_host_w_bits_data, // @[:@25436.4]
  input         io_host_b_ready, // @[:@25436.4]
  output        io_host_b_valid, // @[:@25436.4]
  output        io_host_ar_ready, // @[:@25436.4]
  input         io_host_ar_valid, // @[:@25436.4]
  input  [15:0] io_host_ar_bits_addr, // @[:@25436.4]
  input         io_host_r_ready, // @[:@25436.4]
  output        io_host_r_valid, // @[:@25436.4]
  output [31:0] io_host_r_bits_data, // @[:@25436.4]
  input         io_mem_aw_ready, // @[:@25436.4]
  output        io_mem_aw_valid, // @[:@25436.4]
  output [31:0] io_mem_aw_bits_addr, // @[:@25436.4]
  output [7:0]  io_mem_aw_bits_len, // @[:@25436.4]
  input         io_mem_w_ready, // @[:@25436.4]
  output        io_mem_w_valid, // @[:@25436.4]
  output [63:0] io_mem_w_bits_data, // @[:@25436.4]
  output        io_mem_w_bits_last, // @[:@25436.4]
  output        io_mem_b_ready, // @[:@25436.4]
  input         io_mem_b_valid, // @[:@25436.4]
  input         io_mem_ar_ready, // @[:@25436.4]
  output        io_mem_ar_valid, // @[:@25436.4]
  output [31:0] io_mem_ar_bits_addr, // @[:@25436.4]
  output [7:0]  io_mem_ar_bits_len, // @[:@25436.4]
  output        io_mem_r_ready, // @[:@25436.4]
  input         io_mem_r_valid, // @[:@25436.4]
  input  [63:0] io_mem_r_bits_data, // @[:@25436.4]
  input         io_mem_r_bits_last // @[:@25436.4]
);
  wire  vcr_clock; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_reset; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_aw_ready; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_aw_valid; // @[VTAShell.scala 48:19:@25438.4]
  wire [15:0] vcr_io_host_aw_bits_addr; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_w_ready; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_w_valid; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_host_w_bits_data; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_b_ready; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_b_valid; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_ar_ready; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_ar_valid; // @[VTAShell.scala 48:19:@25438.4]
  wire [15:0] vcr_io_host_ar_bits_addr; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_r_ready; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_host_r_valid; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_host_r_bits_data; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_vcr_launch; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_vcr_finish; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_vcr_ecnt_0_valid; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_vcr_ecnt_0_bits; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_vcr_vals_0; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_vcr_ptrs_0; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_vcr_ptrs_1; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_vcr_ptrs_2; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_vcr_ptrs_3; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_vcr_ptrs_4; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_vcr_ptrs_5; // @[VTAShell.scala 48:19:@25438.4]
  wire  vcr_io_vcr_ucnt_0_valid; // @[VTAShell.scala 48:19:@25438.4]
  wire [31:0] vcr_io_vcr_ucnt_0_bits; // @[VTAShell.scala 48:19:@25438.4]
  wire  vme_clock; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_reset; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_aw_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_aw_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [31:0] vme_io_mem_aw_bits_addr; // @[VTAShell.scala 49:19:@25441.4]
  wire [7:0] vme_io_mem_aw_bits_len; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_w_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_w_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [63:0] vme_io_mem_w_bits_data; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_w_bits_last; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_b_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_b_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_ar_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_ar_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [31:0] vme_io_mem_ar_bits_addr; // @[VTAShell.scala 49:19:@25441.4]
  wire [7:0] vme_io_mem_ar_bits_len; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_r_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_r_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [63:0] vme_io_mem_r_bits_data; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_mem_r_bits_last; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_0_cmd_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_0_cmd_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [31:0] vme_io_vme_rd_0_cmd_bits_addr; // @[VTAShell.scala 49:19:@25441.4]
  wire [7:0] vme_io_vme_rd_0_cmd_bits_len; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_0_data_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_0_data_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [63:0] vme_io_vme_rd_0_data_bits; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_1_cmd_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_1_cmd_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [31:0] vme_io_vme_rd_1_cmd_bits_addr; // @[VTAShell.scala 49:19:@25441.4]
  wire [7:0] vme_io_vme_rd_1_cmd_bits_len; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_1_data_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_1_data_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [63:0] vme_io_vme_rd_1_data_bits; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_2_cmd_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_2_cmd_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [31:0] vme_io_vme_rd_2_cmd_bits_addr; // @[VTAShell.scala 49:19:@25441.4]
  wire [7:0] vme_io_vme_rd_2_cmd_bits_len; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_2_data_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_2_data_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [63:0] vme_io_vme_rd_2_data_bits; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_3_cmd_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_3_cmd_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [31:0] vme_io_vme_rd_3_cmd_bits_addr; // @[VTAShell.scala 49:19:@25441.4]
  wire [7:0] vme_io_vme_rd_3_cmd_bits_len; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_3_data_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_3_data_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [63:0] vme_io_vme_rd_3_data_bits; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_4_cmd_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_4_cmd_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [31:0] vme_io_vme_rd_4_cmd_bits_addr; // @[VTAShell.scala 49:19:@25441.4]
  wire [7:0] vme_io_vme_rd_4_cmd_bits_len; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_4_data_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_rd_4_data_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [63:0] vme_io_vme_rd_4_data_bits; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_wr_0_cmd_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_wr_0_cmd_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [31:0] vme_io_vme_wr_0_cmd_bits_addr; // @[VTAShell.scala 49:19:@25441.4]
  wire [7:0] vme_io_vme_wr_0_cmd_bits_len; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_wr_0_data_ready; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_wr_0_data_valid; // @[VTAShell.scala 49:19:@25441.4]
  wire [63:0] vme_io_vme_wr_0_data_bits; // @[VTAShell.scala 49:19:@25441.4]
  wire  vme_io_vme_wr_0_ack; // @[VTAShell.scala 49:19:@25441.4]
  wire  core_clock; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_reset; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vcr_launch; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vcr_finish; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vcr_ecnt_0_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vcr_ecnt_0_bits; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vcr_vals_0; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vcr_ptrs_0; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vcr_ptrs_1; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vcr_ptrs_2; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vcr_ptrs_3; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vcr_ptrs_4; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vcr_ptrs_5; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vcr_ucnt_0_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vcr_ucnt_0_bits; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_0_cmd_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_0_cmd_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vme_rd_0_cmd_bits_addr; // @[VTAShell.scala 50:20:@25444.4]
  wire [7:0] core_io_vme_rd_0_cmd_bits_len; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_0_data_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_0_data_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [63:0] core_io_vme_rd_0_data_bits; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_1_cmd_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_1_cmd_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vme_rd_1_cmd_bits_addr; // @[VTAShell.scala 50:20:@25444.4]
  wire [7:0] core_io_vme_rd_1_cmd_bits_len; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_1_data_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_1_data_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [63:0] core_io_vme_rd_1_data_bits; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_2_cmd_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_2_cmd_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vme_rd_2_cmd_bits_addr; // @[VTAShell.scala 50:20:@25444.4]
  wire [7:0] core_io_vme_rd_2_cmd_bits_len; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_2_data_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_2_data_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [63:0] core_io_vme_rd_2_data_bits; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_3_cmd_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_3_cmd_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vme_rd_3_cmd_bits_addr; // @[VTAShell.scala 50:20:@25444.4]
  wire [7:0] core_io_vme_rd_3_cmd_bits_len; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_3_data_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_3_data_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [63:0] core_io_vme_rd_3_data_bits; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_4_cmd_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_4_cmd_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vme_rd_4_cmd_bits_addr; // @[VTAShell.scala 50:20:@25444.4]
  wire [7:0] core_io_vme_rd_4_cmd_bits_len; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_4_data_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_rd_4_data_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [63:0] core_io_vme_rd_4_data_bits; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_wr_0_cmd_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_wr_0_cmd_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [31:0] core_io_vme_wr_0_cmd_bits_addr; // @[VTAShell.scala 50:20:@25444.4]
  wire [7:0] core_io_vme_wr_0_cmd_bits_len; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_wr_0_data_ready; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_wr_0_data_valid; // @[VTAShell.scala 50:20:@25444.4]
  wire [63:0] core_io_vme_wr_0_data_bits; // @[VTAShell.scala 50:20:@25444.4]
  wire  core_io_vme_wr_0_ack; // @[VTAShell.scala 50:20:@25444.4]
  VCR vcr ( // @[VTAShell.scala 48:19:@25438.4]
    .clock(vcr_clock),
    .reset(vcr_reset),
    .io_host_aw_ready(vcr_io_host_aw_ready),
    .io_host_aw_valid(vcr_io_host_aw_valid),
    .io_host_aw_bits_addr(vcr_io_host_aw_bits_addr),
    .io_host_w_ready(vcr_io_host_w_ready),
    .io_host_w_valid(vcr_io_host_w_valid),
    .io_host_w_bits_data(vcr_io_host_w_bits_data),
    .io_host_b_ready(vcr_io_host_b_ready),
    .io_host_b_valid(vcr_io_host_b_valid),
    .io_host_ar_ready(vcr_io_host_ar_ready),
    .io_host_ar_valid(vcr_io_host_ar_valid),
    .io_host_ar_bits_addr(vcr_io_host_ar_bits_addr),
    .io_host_r_ready(vcr_io_host_r_ready),
    .io_host_r_valid(vcr_io_host_r_valid),
    .io_host_r_bits_data(vcr_io_host_r_bits_data),
    .io_vcr_launch(vcr_io_vcr_launch),
    .io_vcr_finish(vcr_io_vcr_finish),
    .io_vcr_ecnt_0_valid(vcr_io_vcr_ecnt_0_valid),
    .io_vcr_ecnt_0_bits(vcr_io_vcr_ecnt_0_bits),
    .io_vcr_vals_0(vcr_io_vcr_vals_0),
    .io_vcr_ptrs_0(vcr_io_vcr_ptrs_0),
    .io_vcr_ptrs_1(vcr_io_vcr_ptrs_1),
    .io_vcr_ptrs_2(vcr_io_vcr_ptrs_2),
    .io_vcr_ptrs_3(vcr_io_vcr_ptrs_3),
    .io_vcr_ptrs_4(vcr_io_vcr_ptrs_4),
    .io_vcr_ptrs_5(vcr_io_vcr_ptrs_5),
    .io_vcr_ucnt_0_valid(vcr_io_vcr_ucnt_0_valid),
    .io_vcr_ucnt_0_bits(vcr_io_vcr_ucnt_0_bits)
  );
  VME vme ( // @[VTAShell.scala 49:19:@25441.4]
    .clock(vme_clock),
    .reset(vme_reset),
    .io_mem_aw_ready(vme_io_mem_aw_ready),
    .io_mem_aw_valid(vme_io_mem_aw_valid),
    .io_mem_aw_bits_addr(vme_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(vme_io_mem_aw_bits_len),
    .io_mem_w_ready(vme_io_mem_w_ready),
    .io_mem_w_valid(vme_io_mem_w_valid),
    .io_mem_w_bits_data(vme_io_mem_w_bits_data),
    .io_mem_w_bits_last(vme_io_mem_w_bits_last),
    .io_mem_b_ready(vme_io_mem_b_ready),
    .io_mem_b_valid(vme_io_mem_b_valid),
    .io_mem_ar_ready(vme_io_mem_ar_ready),
    .io_mem_ar_valid(vme_io_mem_ar_valid),
    .io_mem_ar_bits_addr(vme_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(vme_io_mem_ar_bits_len),
    .io_mem_r_ready(vme_io_mem_r_ready),
    .io_mem_r_valid(vme_io_mem_r_valid),
    .io_mem_r_bits_data(vme_io_mem_r_bits_data),
    .io_mem_r_bits_last(vme_io_mem_r_bits_last),
    .io_vme_rd_0_cmd_ready(vme_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(vme_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(vme_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(vme_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(vme_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(vme_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits(vme_io_vme_rd_0_data_bits),
    .io_vme_rd_1_cmd_ready(vme_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(vme_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(vme_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(vme_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_data_ready(vme_io_vme_rd_1_data_ready),
    .io_vme_rd_1_data_valid(vme_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits(vme_io_vme_rd_1_data_bits),
    .io_vme_rd_2_cmd_ready(vme_io_vme_rd_2_cmd_ready),
    .io_vme_rd_2_cmd_valid(vme_io_vme_rd_2_cmd_valid),
    .io_vme_rd_2_cmd_bits_addr(vme_io_vme_rd_2_cmd_bits_addr),
    .io_vme_rd_2_cmd_bits_len(vme_io_vme_rd_2_cmd_bits_len),
    .io_vme_rd_2_data_ready(vme_io_vme_rd_2_data_ready),
    .io_vme_rd_2_data_valid(vme_io_vme_rd_2_data_valid),
    .io_vme_rd_2_data_bits(vme_io_vme_rd_2_data_bits),
    .io_vme_rd_3_cmd_ready(vme_io_vme_rd_3_cmd_ready),
    .io_vme_rd_3_cmd_valid(vme_io_vme_rd_3_cmd_valid),
    .io_vme_rd_3_cmd_bits_addr(vme_io_vme_rd_3_cmd_bits_addr),
    .io_vme_rd_3_cmd_bits_len(vme_io_vme_rd_3_cmd_bits_len),
    .io_vme_rd_3_data_ready(vme_io_vme_rd_3_data_ready),
    .io_vme_rd_3_data_valid(vme_io_vme_rd_3_data_valid),
    .io_vme_rd_3_data_bits(vme_io_vme_rd_3_data_bits),
    .io_vme_rd_4_cmd_ready(vme_io_vme_rd_4_cmd_ready),
    .io_vme_rd_4_cmd_valid(vme_io_vme_rd_4_cmd_valid),
    .io_vme_rd_4_cmd_bits_addr(vme_io_vme_rd_4_cmd_bits_addr),
    .io_vme_rd_4_cmd_bits_len(vme_io_vme_rd_4_cmd_bits_len),
    .io_vme_rd_4_data_ready(vme_io_vme_rd_4_data_ready),
    .io_vme_rd_4_data_valid(vme_io_vme_rd_4_data_valid),
    .io_vme_rd_4_data_bits(vme_io_vme_rd_4_data_bits),
    .io_vme_wr_0_cmd_ready(vme_io_vme_wr_0_cmd_ready),
    .io_vme_wr_0_cmd_valid(vme_io_vme_wr_0_cmd_valid),
    .io_vme_wr_0_cmd_bits_addr(vme_io_vme_wr_0_cmd_bits_addr),
    .io_vme_wr_0_cmd_bits_len(vme_io_vme_wr_0_cmd_bits_len),
    .io_vme_wr_0_data_ready(vme_io_vme_wr_0_data_ready),
    .io_vme_wr_0_data_valid(vme_io_vme_wr_0_data_valid),
    .io_vme_wr_0_data_bits(vme_io_vme_wr_0_data_bits),
    .io_vme_wr_0_ack(vme_io_vme_wr_0_ack)
  );
  Core core ( // @[VTAShell.scala 50:20:@25444.4]
    .clock(core_clock),
    .reset(core_reset),
    .io_vcr_launch(core_io_vcr_launch),
    .io_vcr_finish(core_io_vcr_finish),
    .io_vcr_ecnt_0_valid(core_io_vcr_ecnt_0_valid),
    .io_vcr_ecnt_0_bits(core_io_vcr_ecnt_0_bits),
    .io_vcr_vals_0(core_io_vcr_vals_0),
    .io_vcr_ptrs_0(core_io_vcr_ptrs_0),
    .io_vcr_ptrs_1(core_io_vcr_ptrs_1),
    .io_vcr_ptrs_2(core_io_vcr_ptrs_2),
    .io_vcr_ptrs_3(core_io_vcr_ptrs_3),
    .io_vcr_ptrs_4(core_io_vcr_ptrs_4),
    .io_vcr_ptrs_5(core_io_vcr_ptrs_5),
    .io_vcr_ucnt_0_valid(core_io_vcr_ucnt_0_valid),
    .io_vcr_ucnt_0_bits(core_io_vcr_ucnt_0_bits),
    .io_vme_rd_0_cmd_ready(core_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(core_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(core_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(core_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(core_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(core_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits(core_io_vme_rd_0_data_bits),
    .io_vme_rd_1_cmd_ready(core_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(core_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(core_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(core_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_data_ready(core_io_vme_rd_1_data_ready),
    .io_vme_rd_1_data_valid(core_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits(core_io_vme_rd_1_data_bits),
    .io_vme_rd_2_cmd_ready(core_io_vme_rd_2_cmd_ready),
    .io_vme_rd_2_cmd_valid(core_io_vme_rd_2_cmd_valid),
    .io_vme_rd_2_cmd_bits_addr(core_io_vme_rd_2_cmd_bits_addr),
    .io_vme_rd_2_cmd_bits_len(core_io_vme_rd_2_cmd_bits_len),
    .io_vme_rd_2_data_ready(core_io_vme_rd_2_data_ready),
    .io_vme_rd_2_data_valid(core_io_vme_rd_2_data_valid),
    .io_vme_rd_2_data_bits(core_io_vme_rd_2_data_bits),
    .io_vme_rd_3_cmd_ready(core_io_vme_rd_3_cmd_ready),
    .io_vme_rd_3_cmd_valid(core_io_vme_rd_3_cmd_valid),
    .io_vme_rd_3_cmd_bits_addr(core_io_vme_rd_3_cmd_bits_addr),
    .io_vme_rd_3_cmd_bits_len(core_io_vme_rd_3_cmd_bits_len),
    .io_vme_rd_3_data_ready(core_io_vme_rd_3_data_ready),
    .io_vme_rd_3_data_valid(core_io_vme_rd_3_data_valid),
    .io_vme_rd_3_data_bits(core_io_vme_rd_3_data_bits),
    .io_vme_rd_4_cmd_ready(core_io_vme_rd_4_cmd_ready),
    .io_vme_rd_4_cmd_valid(core_io_vme_rd_4_cmd_valid),
    .io_vme_rd_4_cmd_bits_addr(core_io_vme_rd_4_cmd_bits_addr),
    .io_vme_rd_4_cmd_bits_len(core_io_vme_rd_4_cmd_bits_len),
    .io_vme_rd_4_data_ready(core_io_vme_rd_4_data_ready),
    .io_vme_rd_4_data_valid(core_io_vme_rd_4_data_valid),
    .io_vme_rd_4_data_bits(core_io_vme_rd_4_data_bits),
    .io_vme_wr_0_cmd_ready(core_io_vme_wr_0_cmd_ready),
    .io_vme_wr_0_cmd_valid(core_io_vme_wr_0_cmd_valid),
    .io_vme_wr_0_cmd_bits_addr(core_io_vme_wr_0_cmd_bits_addr),
    .io_vme_wr_0_cmd_bits_len(core_io_vme_wr_0_cmd_bits_len),
    .io_vme_wr_0_data_ready(core_io_vme_wr_0_data_ready),
    .io_vme_wr_0_data_valid(core_io_vme_wr_0_data_valid),
    .io_vme_wr_0_data_bits(core_io_vme_wr_0_data_bits),
    .io_vme_wr_0_ack(core_io_vme_wr_0_ack)
  );
  assign io_host_aw_ready = vcr_io_host_aw_ready; // @[VTAShell.scala 55:15:@25519.4]
  assign io_host_w_ready = vcr_io_host_w_ready; // @[VTAShell.scala 55:15:@25516.4]
  assign io_host_b_valid = vcr_io_host_b_valid; // @[VTAShell.scala 55:15:@25511.4]
  assign io_host_ar_ready = vcr_io_host_ar_ready; // @[VTAShell.scala 55:15:@25509.4]
  assign io_host_r_valid = vcr_io_host_r_valid; // @[VTAShell.scala 55:15:@25505.4]
  assign io_host_r_bits_data = vcr_io_host_r_bits_data; // @[VTAShell.scala 55:15:@25504.4]
  assign io_mem_aw_valid = vme_io_mem_aw_valid; // @[VTAShell.scala 56:10:@25563.4]
  assign io_mem_aw_bits_addr = vme_io_mem_aw_bits_addr; // @[VTAShell.scala 56:10:@25562.4]
  assign io_mem_aw_bits_len = vme_io_mem_aw_bits_len; // @[VTAShell.scala 56:10:@25559.4]
  assign io_mem_w_valid = vme_io_mem_w_valid; // @[VTAShell.scala 56:10:@25550.4]
  assign io_mem_w_bits_data = vme_io_mem_w_bits_data; // @[VTAShell.scala 56:10:@25549.4]
  assign io_mem_w_bits_last = vme_io_mem_w_bits_last; // @[VTAShell.scala 56:10:@25547.4]
  assign io_mem_b_ready = vme_io_mem_b_ready; // @[VTAShell.scala 56:10:@25544.4]
  assign io_mem_ar_valid = vme_io_mem_ar_valid; // @[VTAShell.scala 56:10:@25538.4]
  assign io_mem_ar_bits_addr = vme_io_mem_ar_bits_addr; // @[VTAShell.scala 56:10:@25537.4]
  assign io_mem_ar_bits_len = vme_io_mem_ar_bits_len; // @[VTAShell.scala 56:10:@25534.4]
  assign io_mem_r_ready = vme_io_mem_r_ready; // @[VTAShell.scala 56:10:@25526.4]
  assign vcr_clock = clock; // @[:@25439.4]
  assign vcr_reset = reset; // @[:@25440.4]
  assign vcr_io_host_aw_valid = io_host_aw_valid; // @[VTAShell.scala 55:15:@25518.4]
  assign vcr_io_host_aw_bits_addr = io_host_aw_bits_addr; // @[VTAShell.scala 55:15:@25517.4]
  assign vcr_io_host_w_valid = io_host_w_valid; // @[VTAShell.scala 55:15:@25515.4]
  assign vcr_io_host_w_bits_data = io_host_w_bits_data; // @[VTAShell.scala 55:15:@25514.4]
  assign vcr_io_host_b_ready = io_host_b_ready; // @[VTAShell.scala 55:15:@25512.4]
  assign vcr_io_host_ar_valid = io_host_ar_valid; // @[VTAShell.scala 55:15:@25508.4]
  assign vcr_io_host_ar_bits_addr = io_host_ar_bits_addr; // @[VTAShell.scala 55:15:@25507.4]
  assign vcr_io_host_r_ready = io_host_r_ready; // @[VTAShell.scala 55:15:@25506.4]
  assign vcr_io_vcr_finish = core_io_vcr_finish; // @[VTAShell.scala 52:15:@25458.4]
  assign vcr_io_vcr_ecnt_0_valid = core_io_vcr_ecnt_0_valid; // @[VTAShell.scala 52:15:@25457.4]
  assign vcr_io_vcr_ecnt_0_bits = core_io_vcr_ecnt_0_bits; // @[VTAShell.scala 52:15:@25456.4]
  assign vcr_io_vcr_ucnt_0_valid = core_io_vcr_ucnt_0_valid; // @[VTAShell.scala 52:15:@25448.4]
  assign vcr_io_vcr_ucnt_0_bits = core_io_vcr_ucnt_0_bits; // @[VTAShell.scala 52:15:@25447.4]
  assign vme_clock = clock; // @[:@25442.4]
  assign vme_reset = reset; // @[:@25443.4]
  assign vme_io_mem_aw_ready = io_mem_aw_ready; // @[VTAShell.scala 56:10:@25564.4]
  assign vme_io_mem_w_ready = io_mem_w_ready; // @[VTAShell.scala 56:10:@25551.4]
  assign vme_io_mem_b_valid = io_mem_b_valid; // @[VTAShell.scala 56:10:@25543.4]
  assign vme_io_mem_ar_ready = io_mem_ar_ready; // @[VTAShell.scala 56:10:@25539.4]
  assign vme_io_mem_r_valid = io_mem_r_valid; // @[VTAShell.scala 56:10:@25525.4]
  assign vme_io_mem_r_bits_data = io_mem_r_bits_data; // @[VTAShell.scala 56:10:@25524.4]
  assign vme_io_mem_r_bits_last = io_mem_r_bits_last; // @[VTAShell.scala 56:10:@25522.4]
  assign vme_io_vme_rd_0_cmd_valid = core_io_vme_rd_0_cmd_valid; // @[VTAShell.scala 53:14:@25473.4]
  assign vme_io_vme_rd_0_cmd_bits_addr = core_io_vme_rd_0_cmd_bits_addr; // @[VTAShell.scala 53:14:@25472.4]
  assign vme_io_vme_rd_0_cmd_bits_len = core_io_vme_rd_0_cmd_bits_len; // @[VTAShell.scala 53:14:@25471.4]
  assign vme_io_vme_rd_0_data_ready = core_io_vme_rd_0_data_ready; // @[VTAShell.scala 53:14:@25470.4]
  assign vme_io_vme_rd_1_cmd_valid = core_io_vme_rd_1_cmd_valid; // @[VTAShell.scala 53:14:@25480.4]
  assign vme_io_vme_rd_1_cmd_bits_addr = core_io_vme_rd_1_cmd_bits_addr; // @[VTAShell.scala 53:14:@25479.4]
  assign vme_io_vme_rd_1_cmd_bits_len = core_io_vme_rd_1_cmd_bits_len; // @[VTAShell.scala 53:14:@25478.4]
  assign vme_io_vme_rd_1_data_ready = core_io_vme_rd_1_data_ready; // @[VTAShell.scala 53:14:@25477.4]
  assign vme_io_vme_rd_2_cmd_valid = core_io_vme_rd_2_cmd_valid; // @[VTAShell.scala 53:14:@25487.4]
  assign vme_io_vme_rd_2_cmd_bits_addr = core_io_vme_rd_2_cmd_bits_addr; // @[VTAShell.scala 53:14:@25486.4]
  assign vme_io_vme_rd_2_cmd_bits_len = core_io_vme_rd_2_cmd_bits_len; // @[VTAShell.scala 53:14:@25485.4]
  assign vme_io_vme_rd_2_data_ready = core_io_vme_rd_2_data_ready; // @[VTAShell.scala 53:14:@25484.4]
  assign vme_io_vme_rd_3_cmd_valid = core_io_vme_rd_3_cmd_valid; // @[VTAShell.scala 53:14:@25494.4]
  assign vme_io_vme_rd_3_cmd_bits_addr = core_io_vme_rd_3_cmd_bits_addr; // @[VTAShell.scala 53:14:@25493.4]
  assign vme_io_vme_rd_3_cmd_bits_len = core_io_vme_rd_3_cmd_bits_len; // @[VTAShell.scala 53:14:@25492.4]
  assign vme_io_vme_rd_3_data_ready = core_io_vme_rd_3_data_ready; // @[VTAShell.scala 53:14:@25491.4]
  assign vme_io_vme_rd_4_cmd_valid = core_io_vme_rd_4_cmd_valid; // @[VTAShell.scala 53:14:@25501.4]
  assign vme_io_vme_rd_4_cmd_bits_addr = core_io_vme_rd_4_cmd_bits_addr; // @[VTAShell.scala 53:14:@25500.4]
  assign vme_io_vme_rd_4_cmd_bits_len = core_io_vme_rd_4_cmd_bits_len; // @[VTAShell.scala 53:14:@25499.4]
  assign vme_io_vme_rd_4_data_ready = core_io_vme_rd_4_data_ready; // @[VTAShell.scala 53:14:@25498.4]
  assign vme_io_vme_wr_0_cmd_valid = core_io_vme_wr_0_cmd_valid; // @[VTAShell.scala 53:14:@25466.4]
  assign vme_io_vme_wr_0_cmd_bits_addr = core_io_vme_wr_0_cmd_bits_addr; // @[VTAShell.scala 53:14:@25465.4]
  assign vme_io_vme_wr_0_cmd_bits_len = core_io_vme_wr_0_cmd_bits_len; // @[VTAShell.scala 53:14:@25464.4]
  assign vme_io_vme_wr_0_data_valid = core_io_vme_wr_0_data_valid; // @[VTAShell.scala 53:14:@25462.4]
  assign vme_io_vme_wr_0_data_bits = core_io_vme_wr_0_data_bits; // @[VTAShell.scala 53:14:@25461.4]
  assign core_clock = clock; // @[:@25445.4]
  assign core_reset = reset; // @[:@25446.4]
  assign core_io_vcr_launch = vcr_io_vcr_launch; // @[VTAShell.scala 52:15:@25459.4]
  assign core_io_vcr_vals_0 = vcr_io_vcr_vals_0; // @[VTAShell.scala 52:15:@25455.4]
  assign core_io_vcr_ptrs_0 = vcr_io_vcr_ptrs_0; // @[VTAShell.scala 52:15:@25449.4]
  assign core_io_vcr_ptrs_1 = vcr_io_vcr_ptrs_1; // @[VTAShell.scala 52:15:@25450.4]
  assign core_io_vcr_ptrs_2 = vcr_io_vcr_ptrs_2; // @[VTAShell.scala 52:15:@25451.4]
  assign core_io_vcr_ptrs_3 = vcr_io_vcr_ptrs_3; // @[VTAShell.scala 52:15:@25452.4]
  assign core_io_vcr_ptrs_4 = vcr_io_vcr_ptrs_4; // @[VTAShell.scala 52:15:@25453.4]
  assign core_io_vcr_ptrs_5 = vcr_io_vcr_ptrs_5; // @[VTAShell.scala 52:15:@25454.4]
  assign core_io_vme_rd_0_cmd_ready = vme_io_vme_rd_0_cmd_ready; // @[VTAShell.scala 53:14:@25474.4]
  assign core_io_vme_rd_0_data_valid = vme_io_vme_rd_0_data_valid; // @[VTAShell.scala 53:14:@25469.4]
  assign core_io_vme_rd_0_data_bits = vme_io_vme_rd_0_data_bits; // @[VTAShell.scala 53:14:@25468.4]
  assign core_io_vme_rd_1_cmd_ready = vme_io_vme_rd_1_cmd_ready; // @[VTAShell.scala 53:14:@25481.4]
  assign core_io_vme_rd_1_data_valid = vme_io_vme_rd_1_data_valid; // @[VTAShell.scala 53:14:@25476.4]
  assign core_io_vme_rd_1_data_bits = vme_io_vme_rd_1_data_bits; // @[VTAShell.scala 53:14:@25475.4]
  assign core_io_vme_rd_2_cmd_ready = vme_io_vme_rd_2_cmd_ready; // @[VTAShell.scala 53:14:@25488.4]
  assign core_io_vme_rd_2_data_valid = vme_io_vme_rd_2_data_valid; // @[VTAShell.scala 53:14:@25483.4]
  assign core_io_vme_rd_2_data_bits = vme_io_vme_rd_2_data_bits; // @[VTAShell.scala 53:14:@25482.4]
  assign core_io_vme_rd_3_cmd_ready = vme_io_vme_rd_3_cmd_ready; // @[VTAShell.scala 53:14:@25495.4]
  assign core_io_vme_rd_3_data_valid = vme_io_vme_rd_3_data_valid; // @[VTAShell.scala 53:14:@25490.4]
  assign core_io_vme_rd_3_data_bits = vme_io_vme_rd_3_data_bits; // @[VTAShell.scala 53:14:@25489.4]
  assign core_io_vme_rd_4_cmd_ready = vme_io_vme_rd_4_cmd_ready; // @[VTAShell.scala 53:14:@25502.4]
  assign core_io_vme_rd_4_data_valid = vme_io_vme_rd_4_data_valid; // @[VTAShell.scala 53:14:@25497.4]
  assign core_io_vme_rd_4_data_bits = vme_io_vme_rd_4_data_bits; // @[VTAShell.scala 53:14:@25496.4]
  assign core_io_vme_wr_0_cmd_ready = vme_io_vme_wr_0_cmd_ready; // @[VTAShell.scala 53:14:@25467.4]
  assign core_io_vme_wr_0_data_ready = vme_io_vme_wr_0_data_ready; // @[VTAShell.scala 53:14:@25463.4]
  assign core_io_vme_wr_0_ack = vme_io_vme_wr_0_ack; // @[VTAShell.scala 53:14:@25460.4]
endmodule
module Test( // @[:@25566.2]
  input   clock, // @[:@25567.4]
  input   reset, // @[:@25568.4]
  input   sim_clock, // @[:@25569.4]
  output  sim_wait // @[:@25570.4]
);
  wire  sim_shell_clock; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_reset; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_aw_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_aw_valid; // @[Test.scala 31:25:@25572.4]
  wire [31:0] sim_shell_mem_aw_bits_addr; // @[Test.scala 31:25:@25572.4]
  wire [7:0] sim_shell_mem_aw_bits_len; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_w_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_w_valid; // @[Test.scala 31:25:@25572.4]
  wire [63:0] sim_shell_mem_w_bits_data; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_w_bits_last; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_b_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_b_valid; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_ar_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_ar_valid; // @[Test.scala 31:25:@25572.4]
  wire [31:0] sim_shell_mem_ar_bits_addr; // @[Test.scala 31:25:@25572.4]
  wire [7:0] sim_shell_mem_ar_bits_len; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_r_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_r_valid; // @[Test.scala 31:25:@25572.4]
  wire [63:0] sim_shell_mem_r_bits_data; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_mem_r_bits_last; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_aw_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_aw_valid; // @[Test.scala 31:25:@25572.4]
  wire [15:0] sim_shell_host_aw_bits_addr; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_w_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_w_valid; // @[Test.scala 31:25:@25572.4]
  wire [31:0] sim_shell_host_w_bits_data; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_b_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_b_valid; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_ar_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_ar_valid; // @[Test.scala 31:25:@25572.4]
  wire [15:0] sim_shell_host_ar_bits_addr; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_r_ready; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_host_r_valid; // @[Test.scala 31:25:@25572.4]
  wire [31:0] sim_shell_host_r_bits_data; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_sim_clock; // @[Test.scala 31:25:@25572.4]
  wire  sim_shell_sim_wait; // @[Test.scala 31:25:@25572.4]
  wire  vta_shell_clock; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_reset; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_aw_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_aw_valid; // @[Test.scala 32:25:@25575.4]
  wire [15:0] vta_shell_io_host_aw_bits_addr; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_w_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_w_valid; // @[Test.scala 32:25:@25575.4]
  wire [31:0] vta_shell_io_host_w_bits_data; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_b_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_b_valid; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_ar_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_ar_valid; // @[Test.scala 32:25:@25575.4]
  wire [15:0] vta_shell_io_host_ar_bits_addr; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_r_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_host_r_valid; // @[Test.scala 32:25:@25575.4]
  wire [31:0] vta_shell_io_host_r_bits_data; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_aw_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_aw_valid; // @[Test.scala 32:25:@25575.4]
  wire [31:0] vta_shell_io_mem_aw_bits_addr; // @[Test.scala 32:25:@25575.4]
  wire [7:0] vta_shell_io_mem_aw_bits_len; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_w_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_w_valid; // @[Test.scala 32:25:@25575.4]
  wire [63:0] vta_shell_io_mem_w_bits_data; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_w_bits_last; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_b_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_b_valid; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_ar_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_ar_valid; // @[Test.scala 32:25:@25575.4]
  wire [31:0] vta_shell_io_mem_ar_bits_addr; // @[Test.scala 32:25:@25575.4]
  wire [7:0] vta_shell_io_mem_ar_bits_len; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_r_ready; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_r_valid; // @[Test.scala 32:25:@25575.4]
  wire [63:0] vta_shell_io_mem_r_bits_data; // @[Test.scala 32:25:@25575.4]
  wire  vta_shell_io_mem_r_bits_last; // @[Test.scala 32:25:@25575.4]
  SimShell sim_shell ( // @[Test.scala 31:25:@25572.4]
    .clock(sim_shell_clock),
    .reset(sim_shell_reset),
    .mem_aw_ready(sim_shell_mem_aw_ready),
    .mem_aw_valid(sim_shell_mem_aw_valid),
    .mem_aw_bits_addr(sim_shell_mem_aw_bits_addr),
    .mem_aw_bits_len(sim_shell_mem_aw_bits_len),
    .mem_w_ready(sim_shell_mem_w_ready),
    .mem_w_valid(sim_shell_mem_w_valid),
    .mem_w_bits_data(sim_shell_mem_w_bits_data),
    .mem_w_bits_last(sim_shell_mem_w_bits_last),
    .mem_b_ready(sim_shell_mem_b_ready),
    .mem_b_valid(sim_shell_mem_b_valid),
    .mem_ar_ready(sim_shell_mem_ar_ready),
    .mem_ar_valid(sim_shell_mem_ar_valid),
    .mem_ar_bits_addr(sim_shell_mem_ar_bits_addr),
    .mem_ar_bits_len(sim_shell_mem_ar_bits_len),
    .mem_r_ready(sim_shell_mem_r_ready),
    .mem_r_valid(sim_shell_mem_r_valid),
    .mem_r_bits_data(sim_shell_mem_r_bits_data),
    .mem_r_bits_last(sim_shell_mem_r_bits_last),
    .host_aw_ready(sim_shell_host_aw_ready),
    .host_aw_valid(sim_shell_host_aw_valid),
    .host_aw_bits_addr(sim_shell_host_aw_bits_addr),
    .host_w_ready(sim_shell_host_w_ready),
    .host_w_valid(sim_shell_host_w_valid),
    .host_w_bits_data(sim_shell_host_w_bits_data),
    .host_b_ready(sim_shell_host_b_ready),
    .host_b_valid(sim_shell_host_b_valid),
    .host_ar_ready(sim_shell_host_ar_ready),
    .host_ar_valid(sim_shell_host_ar_valid),
    .host_ar_bits_addr(sim_shell_host_ar_bits_addr),
    .host_r_ready(sim_shell_host_r_ready),
    .host_r_valid(sim_shell_host_r_valid),
    .host_r_bits_data(sim_shell_host_r_bits_data),
    .sim_clock(sim_shell_sim_clock),
    .sim_wait(sim_shell_sim_wait)
  );
  VTAShell vta_shell ( // @[Test.scala 32:25:@25575.4]
    .clock(vta_shell_clock),
    .reset(vta_shell_reset),
    .io_host_aw_ready(vta_shell_io_host_aw_ready),
    .io_host_aw_valid(vta_shell_io_host_aw_valid),
    .io_host_aw_bits_addr(vta_shell_io_host_aw_bits_addr),
    .io_host_w_ready(vta_shell_io_host_w_ready),
    .io_host_w_valid(vta_shell_io_host_w_valid),
    .io_host_w_bits_data(vta_shell_io_host_w_bits_data),
    .io_host_b_ready(vta_shell_io_host_b_ready),
    .io_host_b_valid(vta_shell_io_host_b_valid),
    .io_host_ar_ready(vta_shell_io_host_ar_ready),
    .io_host_ar_valid(vta_shell_io_host_ar_valid),
    .io_host_ar_bits_addr(vta_shell_io_host_ar_bits_addr),
    .io_host_r_ready(vta_shell_io_host_r_ready),
    .io_host_r_valid(vta_shell_io_host_r_valid),
    .io_host_r_bits_data(vta_shell_io_host_r_bits_data),
    .io_mem_aw_ready(vta_shell_io_mem_aw_ready),
    .io_mem_aw_valid(vta_shell_io_mem_aw_valid),
    .io_mem_aw_bits_addr(vta_shell_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(vta_shell_io_mem_aw_bits_len),
    .io_mem_w_ready(vta_shell_io_mem_w_ready),
    .io_mem_w_valid(vta_shell_io_mem_w_valid),
    .io_mem_w_bits_data(vta_shell_io_mem_w_bits_data),
    .io_mem_w_bits_last(vta_shell_io_mem_w_bits_last),
    .io_mem_b_ready(vta_shell_io_mem_b_ready),
    .io_mem_b_valid(vta_shell_io_mem_b_valid),
    .io_mem_ar_ready(vta_shell_io_mem_ar_ready),
    .io_mem_ar_valid(vta_shell_io_mem_ar_valid),
    .io_mem_ar_bits_addr(vta_shell_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(vta_shell_io_mem_ar_bits_len),
    .io_mem_r_ready(vta_shell_io_mem_r_ready),
    .io_mem_r_valid(vta_shell_io_mem_r_valid),
    .io_mem_r_bits_data(vta_shell_io_mem_r_bits_data),
    .io_mem_r_bits_last(vta_shell_io_mem_r_bits_last)
  );
  assign sim_wait = sim_shell_sim_wait; // @[Test.scala 34:12:@25579.4]
  assign sim_shell_clock = clock; // @[:@25573.4]
  assign sim_shell_reset = reset; // @[:@25574.4]
  assign sim_shell_mem_aw_valid = vta_shell_io_mem_aw_valid; // @[Test.scala 35:17:@25623.4]
  assign sim_shell_mem_aw_bits_addr = vta_shell_io_mem_aw_bits_addr; // @[Test.scala 35:17:@25622.4]
  assign sim_shell_mem_aw_bits_len = vta_shell_io_mem_aw_bits_len; // @[Test.scala 35:17:@25619.4]
  assign sim_shell_mem_w_valid = vta_shell_io_mem_w_valid; // @[Test.scala 35:17:@25610.4]
  assign sim_shell_mem_w_bits_data = vta_shell_io_mem_w_bits_data; // @[Test.scala 35:17:@25609.4]
  assign sim_shell_mem_w_bits_last = vta_shell_io_mem_w_bits_last; // @[Test.scala 35:17:@25607.4]
  assign sim_shell_mem_b_ready = vta_shell_io_mem_b_ready; // @[Test.scala 35:17:@25604.4]
  assign sim_shell_mem_ar_valid = vta_shell_io_mem_ar_valid; // @[Test.scala 35:17:@25598.4]
  assign sim_shell_mem_ar_bits_addr = vta_shell_io_mem_ar_bits_addr; // @[Test.scala 35:17:@25597.4]
  assign sim_shell_mem_ar_bits_len = vta_shell_io_mem_ar_bits_len; // @[Test.scala 35:17:@25594.4]
  assign sim_shell_mem_r_ready = vta_shell_io_mem_r_ready; // @[Test.scala 35:17:@25586.4]
  assign sim_shell_host_aw_ready = vta_shell_io_host_aw_ready; // @[Test.scala 36:21:@25641.4]
  assign sim_shell_host_w_ready = vta_shell_io_host_w_ready; // @[Test.scala 36:21:@25638.4]
  assign sim_shell_host_b_valid = vta_shell_io_host_b_valid; // @[Test.scala 36:21:@25633.4]
  assign sim_shell_host_ar_ready = vta_shell_io_host_ar_ready; // @[Test.scala 36:21:@25631.4]
  assign sim_shell_host_r_valid = vta_shell_io_host_r_valid; // @[Test.scala 36:21:@25627.4]
  assign sim_shell_host_r_bits_data = vta_shell_io_host_r_bits_data; // @[Test.scala 36:21:@25626.4]
  assign sim_shell_sim_clock = sim_clock; // @[Test.scala 33:23:@25578.4]
  assign vta_shell_clock = clock; // @[:@25576.4]
  assign vta_shell_reset = reset; // @[:@25577.4]
  assign vta_shell_io_host_aw_valid = sim_shell_host_aw_valid; // @[Test.scala 36:21:@25640.4]
  assign vta_shell_io_host_aw_bits_addr = sim_shell_host_aw_bits_addr; // @[Test.scala 36:21:@25639.4]
  assign vta_shell_io_host_w_valid = sim_shell_host_w_valid; // @[Test.scala 36:21:@25637.4]
  assign vta_shell_io_host_w_bits_data = sim_shell_host_w_bits_data; // @[Test.scala 36:21:@25636.4]
  assign vta_shell_io_host_b_ready = sim_shell_host_b_ready; // @[Test.scala 36:21:@25634.4]
  assign vta_shell_io_host_ar_valid = sim_shell_host_ar_valid; // @[Test.scala 36:21:@25630.4]
  assign vta_shell_io_host_ar_bits_addr = sim_shell_host_ar_bits_addr; // @[Test.scala 36:21:@25629.4]
  assign vta_shell_io_host_r_ready = sim_shell_host_r_ready; // @[Test.scala 36:21:@25628.4]
  assign vta_shell_io_mem_aw_ready = sim_shell_mem_aw_ready; // @[Test.scala 35:17:@25624.4]
  assign vta_shell_io_mem_w_ready = sim_shell_mem_w_ready; // @[Test.scala 35:17:@25611.4]
  assign vta_shell_io_mem_b_valid = sim_shell_mem_b_valid; // @[Test.scala 35:17:@25603.4]
  assign vta_shell_io_mem_ar_ready = sim_shell_mem_ar_ready; // @[Test.scala 35:17:@25599.4]
  assign vta_shell_io_mem_r_valid = sim_shell_mem_r_valid; // @[Test.scala 35:17:@25585.4]
  assign vta_shell_io_mem_r_bits_data = sim_shell_mem_r_bits_data; // @[Test.scala 35:17:@25584.4]
  assign vta_shell_io_mem_r_bits_last = sim_shell_mem_r_bits_last; // @[Test.scala 35:17:@25582.4]
endmodule
